�(]q (cenvironment
an_object
q)�q}q(X   obj_idqKX   positionqcenvironment
position
q)�q}q(X   xq	G?�\(�X   yq
G?�      ubX   colourqX   bqX   shapeqX   circleqX   last_actionqG�      X   current_zoneqKubh)�q}q(hKhh)�q}q(h	G��=p��
=h
G?�333333ubhhhhhG�      hKubh)�q}q(hKhh)�q}q(h	G���
=p��h
G��Q��ubhhhhhG�      hKubh)�q}q(hKhh)�q}q(h	G��G�z�Hh
G?θQ��ubhX   gqhX   triangleqhG�      hKubh)�q}q (hKhh)�q!}q"(h	G��z�G�{h
G?���Q�ubhX   rq#hhhG�      hKubh)�q$}q%(hKhh)�q&}q'(h	G����Q�h
G���\(�ubhhhX   squareq(hG�      hKubh)�q)}q*(hKhh)�q+}q,(h	G?�\(�\h
G?��\(�ubhh#hhhG�      hKubh)�q-}q.(hKhh)�q/}q0(h	G?�\(�h
G��p��
=qubhhhhhG�      hKubh)�q1}q2(hK	hh)�q3}q4(h	G?ۅ�Q�h
G��Q��RubhhhhhG�      hKubh)�q5}q6(hK
hh)�q7}q8(h	G?�G�z�Hh
G��������ubhh#hhhG�      hKubh)�q9}q:(hKhh)�q;}q<(h	G?�G�z�Hh
G��
=p��
ubhhhh(hG�      hKubh)�q=}q>(hKhh)�q?}q@(h	G?�333333h
G��(�\)ubhhhhhG�      hKubh)�qA}qB(hKhh)�qC}qD(h	G?���Q�h
G���Q�ubhh#hhhG�      hKubh)�qE}qF(hKhh)�qG}qH(h	G���G�z�h
G��\(�\ubhhhhhG�      hKubh)�qI}qJ(hKhh)�qK}qL(h	G���
=p�h
G��z�G�{ubhhhhhG�      hKubh)�qM}qN(hKhh)�qO}qP(h	G��(�\)h
G��      ubhhhhhG�      hKubh)�qQ}qR(hKhh)�qS}qT(h	G����Q�h
G?�z�G�ubhhhhhG�      hKubh)�qU}qV(hKhh)�qW}qX(h	G����Q�h
G��\(�ubhhhhhG�      hKubh)�qY}qZ(hKhh)�q[}q\(h	G?�      h
G?��G�z�ubhhhhhG�      hKubh)�q]}q^(hKhh)�q_}q`(h	G?��Q�h
G?�z�G�ubhhhh(hG�      hKubh)�qa}qb(hKhh)�qc}qd(h	G?�333333h
G?�������ubhh#hhhG�      hKubh)�qe}qf(hKhh)�qg}qh(h	G�ٙ�����h
G��z�G�ubhhhhhG�      hKubh)�qi}qj(hKhh)�qk}ql(h	G���Q��h
G����Q�ubhhhh(hG�      hKubh)�qm}qn(hKhh)�qo}qp(h	G�ə�����h
G��\(��ubhhhhhG�      hKubh)�qq}qr(hKhh)�qs}qt(h	G?�Q��h
G��z�G�ubhh#hhhG�      hKubh)�qu}qv(hKhh)�qw}qx(h	G?θQ��h
G��333333ubhh#hhhG�      hKubh)�qy}qz(hKhh)�q{}q|(h	G?�������h
G?陙����ubhhhhhG�      hKubh)�q}}q~(hKhh)�q}q�(h	G?�      h
G���
=p��ubhh#hhhG�      hKubh)�q�}q�(hKhh)�q�}q�(h	G��Q��Rh
G?�333333ubhhhhhG�      hKubh)�q�}q�(hKhh)�q�}q�(h	G?�p��
=qh
G?�\(��ubhh#hhhG�      hKubh)�q�}q�(hKhh)�q�}q�(h	G?�Q��Rh
G?�
=p��
ubhh#hh(hG�      hKubh)�q�}q�(hK hh)�q�}q�(h	G����Q�h
G�У�
=p�ubhh#hhhG�      hKubh)�q�}q�(hK!hh)�q�}q�(h	G?��\(�h
G��p��
=qubhh#hh(hG�      hKubh)�q�}q�(hK"hh)�q�}q�(h	G��p��
=qh
G?�
=p��
ubhh#hhhG�      hKubh)�q�}q�(hK#hh)�q�}q�(h	G��
=p��
h
G��333333ubhh#hhhG�      hKubh)�q�}q�(hK$hh)�q�}q�(h	G��G�z�Hh
G��
=p��
ubhhhhhG�      hKubh)�q�}q�(hK%hh)�q�}q�(h	G��      h
G?�p��
=qubhh#hhhG�      hKubh)�q�}q�(hK&hh)�q�}q�(h	G����Q�h
G��(�\)ubhhhh(hG�      hKubh)�q�}q�(hK'hh)�q�}q�(h	G��ffffffh
G?��G�z�ubhhhhhG�      hKubh)�q�}q�(hK(hh)�q�}q�(h	G?��Q��h
G?��G�z�ubhhhhhG�      hKube]q�(h#hhe]q�(h(hhe}q�(KG��UUUUUVKG?�UUUUUTKG?�      utq�.