�]q (]q(X   Normsq]q(X   Oblq]q(X   Movedq]q(X   ColourqX   anyq	e]q
(X   Shapeqh	e]q(X   ZoneqX   2qe]q(X   Movedq]q(hX   bqe]q(hX   triangleqe]q(hhe]q(X	   Next-Moveq]q(hh	e]q(hX   squareqeeee]q(hhee]q(X   Perq]q(X   ActionqX   putdownq e]q!(hX   gq"e]q#(hhe]q$(X   PerZoneq%X   3q&eeehh]q'(h]q((h]q)(h]q*(hh	e]q+(hh	e]q,(hhe]q-(h]q.(hh	e]q/(hhe]q0(hhe]q1(h]q2(hh	e]q3(hheeee]q4(hhee]q5(h]q6(hh e]q7(hh"e]q8(hhe]q9(h%h&eeeh']q:(h]q;(h]q<(h]q=(hh	e]q>(hh	e]q?(hhe]q@(h]qA(hh	e]qB(hhe]qC(hhe]qD(h]qE(hh	e]qF(hheeee]qG(hhee]qH(h]qI(hh e]qJ(hh"e]qK(hhe]qL(h%h&eeeh:h:h:h:h:h:h:h:h:h:h:h:h:h:h:h:h:h:h:h:h:h:h:h:h:]qM(h]qN(h]qO(h]qP(hh	e]qQ(hh	e]qR(hhe]qS(h]qT(hh	e]qU(hhe]qV(hhe]qW(h]qX(hh	e]qY(hheeee]qZ(hhee]q[(h]q\(hh e]q](hh"e]q^(hhe]q_(h%h&eee]q`(h]qa(h]qb(h]qc(hh	e]qd(hh	e]qe(hhe]qf(h]qg(hh	e]qh(hhe]qi(hhe]qj(h]qk(hh	e]ql(hheeee]qm(hhee]qn(h]qo(hh e]qp(hh"e]qq(hh	e]qr(h%h&eee]qs(h]qt(h]qu(h]qv(hh	e]qw(hh	e]qx(hhe]qy(h]qz(hh	e]q{(hhe]q|(hhe]q}(h]q~(hh	e]q(hheeee]q�(hhee]q�(h]q�(hh e]q�(hh"e]q�(hh	e]q�(h%h&eeehshs]q�(h]q�(h]q�(h]q�(hh	e]q�(hh	e]q�(hhe]q�(h]q�(hh	e]q�(hhe]q�(hhe]q�(h]q�(hh	e]q�(hheeee]q�(hhee]q�(h]q�(hh e]q�(hh"e]q�(hh	e]q�(h%h&eeeh�h�h�]q�(h]q�(h]q�(h]q�(hh	e]q�(hh	e]q�(hhe]q�(h]q�(hh	e]q�(hhe]q�(hhe]q�(h]q�(hh	e]q�(hheeee]q�(hhee]q�(h]q�(hh e]q�(hh"e]q�(hh	e]q�(h%h&eeeh�]q�(h]q�(h]q�(h]q�(hh	e]q�(hh	e]q�(hhe]q�(h]q�(hh	e]q�(hhe]q�(hhe]q�(h]q�(hh	e]q�(hheeee]q�(hhee]q�(h]q�(hh e]q�(hh"e]q�(hh	e]q�(h%h&eee]q�(h]q�(h]q�(h]q�(hh	e]q�(hh	e]q�(hhe]q�(h]q�(hh	e]q�(hhe]q�(hhe]q�(h]q�(hh	e]q�(hheeee]q�(hhee]q�(h]q�(hh e]q�(hh"e]q�(hh	e]q�(h%h&eee]q�(h]q�(h]q�(h]q�(hh	e]q�(hh	e]q�(hhe]q�(h]q�(hh	e]q�(hhe]q�(hhe]q�(h]q�(hh	e]q�(hheeee]q�(hhee]q�(h]q�(hh e]q�(hh"e]q�(hh	e]q�(h%h&eeeh�h�]q�(h]q�(h]q�(h]q�(hh	e]q�(hh	e]q�(hhe]q�(h]q�(hh	e]q�(hhe]q�(hhe]q�(h]q�(hh	e]q�(hheeee]q�(hhee]q�(h]q�(hh e]q�(hh"e]q�(hh	e]q�(h%h&eeeh�h�h�h�]q�(h]q�(h]q�(h]q�(hh	e]q�(hh	e]q�(hhe]q�(h]q�(hh	e]r   (hhe]r  (hhe]r  (h]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r	  (hh	e]r
  (h%h&eee]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hh	e]r  (hhe]r  (hhe]r  (h]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hh	e]r  (h%h&eeej  ]r  (h]r  (h]r   (h]r!  (hh	e]r"  (hh	e]r#  (hhe]r$  (h]r%  (hh	e]r&  (hhe]r'  (hhe]r(  (h]r)  (hh	e]r*  (hheeee]r+  (hhee]r,  (h]r-  (hh e]r.  (hh"e]r/  (hh	e]r0  (h%h&eeej  j  j  ]r1  (h]r2  (h]r3  (h]r4  (hh	e]r5  (hh	e]r6  (hhe]r7  (h]r8  (hh	e]r9  (hhe]r:  (hhe]r;  (h]r<  (hh	e]r=  (hheeee]r>  (hhee]r?  (h]r@  (hh e]rA  (hh"e]rB  (hh	e]rC  (h%h&eeej1  j1  j1  ]rD  (h]rE  (h]rF  (h]rG  (hh	e]rH  (hh	e]rI  (hhe]rJ  (h]rK  (hh	e]rL  (hhe]rM  (hhe]rN  (h]rO  (hh	e]rP  (hheeee]rQ  (hhee]rR  (h]rS  (hh e]rT  (hh"e]rU  (hh	e]rV  (h%h&eeejD  jD  ]rW  (h]rX  (h]rY  (h]rZ  (hh	e]r[  (hh	e]r\  (hhe]r]  (h]r^  (hh	e]r_  (hhe]r`  (hhe]ra  (h]rb  (hh	e]rc  (hheeee]rd  (hhee]re  (h]rf  (hh e]rg  (hh"e]rh  (hh	e]ri  (h%h&eeejW  jW  jW  jW  jW  ]rj  (h]rk  (h]rl  (h]rm  (hh	e]rn  (hh	e]ro  (hhe]rp  (h]rq  (hh	e]rr  (hhe]rs  (hhe]rt  (h]ru  (hh	e]rv  (hheeee]rw  (hhee]rx  (h]ry  (hh e]rz  (hh"e]r{  (hh	e]r|  (h%h&eeejj  ]r}  (h]r~  (h]r  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r   (hhe]r  (h%h&eeej�  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r	  (hh	e]r
  (hhe]r  (hhe]r  (h]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hhe]r  (h%h&eeej  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hh	e]r  (hhe]r  (hhe]r  (h]r   (hh	e]r!  (hheeee]r"  (hhee]r#  (h]r$  (hh e]r%  (hh"e]r&  (hhe]r'  (h%h&eeej  j  j  j  j  ]r(  (h]r)  (h]r*  (h]r+  (hh	e]r,  (hh	e]r-  (hhe]r.  (h]r/  (hh	e]r0  (hhe]r1  (hhe]r2  (h]r3  (hh	e]r4  (hheeee]r5  (hhee]r6  (h]r7  (hh e]r8  (hh"e]r9  (hhe]r:  (h%h&eeej(  j(  j(  j(  j(  j(  j(  j(  j(  j(  j(  j(  ]r;  (h]r<  (h]r=  (h]r>  (hh	e]r?  (hh	e]r@  (hhe]rA  (h]rB  (hh	e]rC  (hhe]rD  (hhe]rE  (h]rF  (hh	e]rG  (hheeee]rH  (hhee]rI  (h]rJ  (hh e]rK  (hh"e]rL  (hhe]rM  (h%h&eeej;  j;  j;  ]rN  (h]rO  (h]rP  (h]rQ  (hh	e]rR  (hh	e]rS  (hhe]rT  (h]rU  (hh	e]rV  (hhe]rW  (hhe]rX  (h]rY  (hh	e]rZ  (hheeee]r[  (hhee]r\  (h]r]  (hh e]r^  (hh"e]r_  (hhe]r`  (h%h&eeejN  ]ra  (h]rb  (h]rc  (h]rd  (hh	e]re  (hh	e]rf  (hhe]rg  (h]rh  (hh	e]ri  (hhe]rj  (hhe]rk  (h]rl  (hh	e]rm  (hheeee]rn  (hhee]ro  (h]rp  (hh e]rq  (hh"e]rr  (hhe]rs  (h%h&eeeja  ja  ja  ]rt  (h]ru  (h]rv  (h]rw  (hh	e]rx  (hh	e]ry  (hhe]rz  (h]r{  (hh	e]r|  (hhe]r}  (hhe]r~  (h]r  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r   (hh	e]r  (hhe]r  (hhe]r  (h]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r	  (hh"e]r
  (hh	e]r  (h%h&eeej�  j�  j�  j�  j�  j�  j�  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hh	e]r  (hhe]r  (hhe]r  (h]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hh	e]r  (h%h&eee]r  (h]r   (h]r!  (h]r"  (hh	e]r#  (hh	e]r$  (hhe]r%  (h]r&  (hh	e]r'  (hhe]r(  (hhe]r)  (h]r*  (hh	e]r+  (hheeee]r,  (hhee]r-  (h]r.  (hh e]r/  (hh"e]r0  (hh	e]r1  (h%h&eeej  j  j  j  ]r2  (h]r3  (h]r4  (h]r5  (hh	e]r6  (hh	e]r7  (hhe]r8  (h]r9  (hh	e]r:  (hhe]r;  (hhe]r<  (h]r=  (hh	e]r>  (hheeee]r?  (hhee]r@  (h]rA  (hh e]rB  (hh"e]rC  (hh	e]rD  (h%h&eeej2  ]rE  (h]rF  (h]rG  (h]rH  (hh	e]rI  (hh	e]rJ  (hhe]rK  (h]rL  (hh	e]rM  (hhe]rN  (hhe]rO  (h]rP  (hh	e]rQ  (hheeee]rR  (hhee]rS  (h]rT  (hh e]rU  (hh"e]rV  (hh	e]rW  (h%h&eee]rX  (h]rY  (h]rZ  (h]r[  (hh	e]r\  (hh	e]r]  (hhe]r^  (h]r_  (hh	e]r`  (hhe]ra  (hhe]rb  (h]rc  (hh	e]rd  (hheeee]re  (hhee]rf  (h]rg  (hh e]rh  (hh"e]ri  (hh	e]rj  (h%h&eeejX  jX  jX  jX  ]rk  (h]rl  (h]rm  (h]rn  (hh	e]ro  (hh	e]rp  (hhe]rq  (h]rr  (hh	e]rs  (hhe]rt  (hhe]ru  (h]rv  (hh	e]rw  (hheeee]rx  (hhee]ry  (h]rz  (hh e]r{  (hh"e]r|  (hh	e]r}  (h%h&eeejk  jk  jk  jk  jk  jk  jk  ]r~  (h]r  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej~  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r   (hh"e]r  (hh	e]r  (h%h&eeej�  j�  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r	  (h]r
  (hh	e]r  (hhe]r  (hhe]r  (h]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hh	e]r  (h%h&eeej  j  j  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hh	e]r  (hhe]r  (hhe]r   (h]r!  (hh	e]r"  (hheeee]r#  (hhee]r$  (h]r%  (hh e]r&  (hh"e]r'  (hh	e]r(  (h%h&eeej  j  j  j  j  j  j  ]r)  (h]r*  (h]r+  (h]r,  (hh	e]r-  (hh	e]r.  (hhe]r/  (h]r0  (hh	e]r1  (hhe]r2  (hhe]r3  (h]r4  (hh	e]r5  (hheeee]r6  (hhee]r7  (h]r8  (hh e]r9  (hh"e]r:  (hhe]r;  (h%h&eeej)  ]r<  (h]r=  (h]r>  (h]r?  (hh	e]r@  (hh	e]rA  (hhe]rB  (h]rC  (hh	e]rD  (hhe]rE  (hhe]rF  (h]rG  (hh	e]rH  (hheeee]rI  (hhee]rJ  (h]rK  (hh e]rL  (hh"e]rM  (hhe]rN  (h%h&eeej<  j<  j<  j<  j<  j<  ]rO  (h]rP  (h]rQ  (h]rR  (hh	e]rS  (hh	e]rT  (hhe]rU  (h]rV  (hh	e]rW  (hhe]rX  (hhe]rY  (h]rZ  (hh	e]r[  (hheeee]r\  (hhee]r]  (h]r^  (hh e]r_  (hh"e]r`  (hhe]ra  (h%h&eeejO  ]rb  (h]rc  (h]rd  (h]re  (hh	e]rf  (hh	e]rg  (hhe]rh  (h]ri  (hh	e]rj  (hhe]rk  (hhe]rl  (h]rm  (hh	e]rn  (hheeee]ro  (hhee]rp  (h]rq  (hh e]rr  (hh"e]rs  (hhe]rt  (h%h&eee]ru  (h]rv  (h]rw  (h]rx  (hh	e]ry  (hh	e]rz  (hhe]r{  (h]r|  (hh	e]r}  (hhe]r~  (hhe]r  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeeju  ju  ju  ju  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r   (h]r  (hhe]r  (hhe]r  (hhe]r  (h]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r	  (hh e]r
  (hh"e]r  (hhe]r  (h%h&eeej�  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r  (hhe]r  (h]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hhe]r  (h%h&eee]r   (h]r!  (h]r"  (h]r#  (hh	e]r$  (hh	e]r%  (hhe]r&  (h]r'  (hhe]r(  (hhe]r)  (hhe]r*  (h]r+  (hh	e]r,  (hheeee]r-  (hhee]r.  (h]r/  (hh e]r0  (hh"e]r1  (hh	e]r2  (h%h&eeej   j   ]r3  (h]r4  (h]r5  (h]r6  (hh	e]r7  (hh	e]r8  (hhe]r9  (h]r:  (hhe]r;  (hhe]r<  (hhe]r=  (h]r>  (hh	e]r?  (hheeee]r@  (hhee]rA  (h]rB  (hh e]rC  (hh"e]rD  (hh	e]rE  (h%h&eeej3  j3  ]rF  (h]rG  (h]rH  (h]rI  (hh	e]rJ  (hh	e]rK  (hhe]rL  (h]rM  (hhe]rN  (hhe]rO  (hhe]rP  (h]rQ  (hh	e]rR  (hheeee]rS  (hhee]rT  (h]rU  (hh e]rV  (hh"e]rW  (hh	e]rX  (h%h&eeejF  jF  jF  jF  jF  jF  ]rY  (h]rZ  (h]r[  (h]r\  (hh	e]r]  (hh	e]r^  (hhe]r_  (h]r`  (hhe]ra  (hhe]rb  (hhe]rc  (h]rd  (hh	e]re  (hheeee]rf  (hhee]rg  (h]rh  (hh e]ri  (hh"e]rj  (hh	e]rk  (h%h&eeejY  jY  jY  jY  jY  ]rl  (h]rm  (h]rn  (h]ro  (hh	e]rp  (hh	e]rq  (hhe]rr  (h]rs  (hhe]rt  (hhe]ru  (hhe]rv  (h]rw  (hh	e]rx  (hheeee]ry  (hhee]rz  (h]r{  (hh e]r|  (hh"e]r}  (hh	e]r~  (h%h&eeejl  jl  jl  jl  ]r  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej  j  j  j  j  j  j  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r   (hh e]r  (hh"e]r  (hh	e]r  (h%h&eeej�  j�  j�  j�  j�  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r	  (hhe]r
  (h]r  (hhe]r  (hhe]r  (hhe]r  (h]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hh	e]r  (h%h&eeej  j  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r   (hhe]r!  (h]r"  (hh	e]r#  (hheeee]r$  (hhee]r%  (h]r&  (hh e]r'  (hh"e]r(  (hh	e]r)  (h%h&eeej  j  ]r*  (h]r+  (h]r,  (h]r-  (hh	e]r.  (hh	e]r/  (hhe]r0  (h]r1  (hhe]r2  (hhe]r3  (hhe]r4  (h]r5  (hh	e]r6  (hheeee]r7  (hhee]r8  (h]r9  (hh e]r:  (hh"e]r;  (hh	e]r<  (h%h&eeej*  j*  ]r=  (h]r>  (h]r?  (h]r@  (hh	e]rA  (hh	e]rB  (hhe]rC  (h]rD  (hhe]rE  (hhe]rF  (hhe]rG  (h]rH  (hh	e]rI  (hheeee]rJ  (hhee]rK  (h]rL  (hh e]rM  (hh"e]rN  (hh	e]rO  (h%h&eee]rP  (h]rQ  (h]rR  (h]rS  (hh	e]rT  (hh	e]rU  (hhe]rV  (h]rW  (hhe]rX  (hhe]rY  (hhe]rZ  (h]r[  (hh	e]r\  (hheeee]r]  (hhee]r^  (h]r_  (hh e]r`  (hh"e]ra  (hh	e]rb  (h%h&eeejP  jP  jP  ]rc  (h]rd  (h]re  (h]rf  (hh	e]rg  (hh	e]rh  (hhe]ri  (h]rj  (hhe]rk  (hhe]rl  (hhe]rm  (h]rn  (hh	e]ro  (hheeee]rp  (hhee]rq  (h]rr  (hh e]rs  (hh"e]rt  (hhe]ru  (h%h&eeejc  jc  jc  jc  jc  jc  jc  jc  ]rv  (h]rw  (h]rx  (h]ry  (hh	e]rz  (hh	e]r{  (hhe]r|  (h]r}  (hhe]r~  (hhe]r  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeejv  jv  jv  jv  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (h]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (X	   Next-Mover�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r   (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r  (hhe]r  (j�  ]r  (hh	e]r  (hheeee]r	  (hhee]r
  (h]r  (hh e]r  (hh"e]r  (hhe]r  (h%h&eeej�  j�  j�  j�  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r  (hhe]r  (j�  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r   (hhe]r!  (h%h&eee]r"  (h]r#  (h]r$  (h]r%  (hh	e]r&  (hh	e]r'  (hhe]r(  (h]r)  (hhe]r*  (hhe]r+  (hhe]r,  (j�  ]r-  (hh	e]r.  (hheeee]r/  (hhee]r0  (h]r1  (hh e]r2  (hh"e]r3  (hhe]r4  (h%h&eeej"  ]r5  (h]r6  (h]r7  (h]r8  (hh	e]r9  (hh	e]r:  (hhe]r;  (h]r<  (hhe]r=  (hhe]r>  (hhe]r?  (j�  ]r@  (hh	e]rA  (hheeee]rB  (hhee]rC  (h]rD  (hh e]rE  (hh"e]rF  (hhe]rG  (h%h&eeej5  j5  j5  ]rH  (h]rI  (h]rJ  (h]rK  (hh	e]rL  (hh	e]rM  (hhe]rN  (h]rO  (hhe]rP  (hhe]rQ  (hhe]rR  (j�  ]rS  (hh	e]rT  (hheeee]rU  (hhee]rV  (h]rW  (hh e]rX  (hh"e]rY  (hhe]rZ  (h%h&eeejH  jH  jH  jH  ]r[  (h]r\  (h]r]  (h]r^  (hh	e]r_  (hh	e]r`  (hhe]ra  (h]rb  (hhe]rc  (hhe]rd  (hhe]re  (j�  ]rf  (hh	e]rg  (hheeee]rh  (hhee]ri  (h]rj  (hh e]rk  (hh"e]rl  (hhe]rm  (h%h&eeej[  j[  ]rn  (h]ro  (h]rp  (h]rq  (hh	e]rr  (hh	e]rs  (hhe]rt  (h]ru  (hhe]rv  (hhe]rw  (hhe]rx  (j�  ]ry  (hh	e]rz  (hheeee]r{  (hhee]r|  (h]r}  (hh e]r~  (hh"e]r  (hhe]r�  (h%h&eeejn  jn  jn  jn  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r   (hhee]r  (h]r  (hh e]r  (hh"e]r  (hhe]r  (h%h&eee]r  (h]r  (h]r  (h]r	  (hh	e]r
  (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r  (hhe]r  (j�  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hhe]r  (h%h&eeej  j  j  j  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r   (hh	e]r!  (hhe]r"  (hhe]r#  (j�  ]r$  (hh	e]r%  (hheeee]r&  (hhee]r'  (h]r(  (hh e]r)  (hh"e]r*  (hhe]r+  (h%h&eeej  j  j  j  j  j  j  ]r,  (h]r-  (h]r.  (h]r/  (hh	e]r0  (hh	e]r1  (hhe]r2  (h]r3  (hh	e]r4  (hhe]r5  (hhe]r6  (j�  ]r7  (hh	e]r8  (hheeee]r9  (hhee]r:  (h]r;  (hh e]r<  (hh"e]r=  (hhe]r>  (h%h&eee]r?  (h]r@  (h]rA  (h]rB  (hh	e]rC  (hh	e]rD  (hhe]rE  (h]rF  (hh	e]rG  (hhe]rH  (hhe]rI  (j�  ]rJ  (hh	e]rK  (hheeee]rL  (hhee]rM  (h]rN  (hh e]rO  (hh"e]rP  (hhe]rQ  (h%h&eeej?  j?  ]rR  (h]rS  (h]rT  (h]rU  (hh	e]rV  (hh	e]rW  (hhe]rX  (h]rY  (hh	e]rZ  (hhe]r[  (hhe]r\  (j�  ]r]  (hh	e]r^  (hheeee]r_  (hhee]r`  (h]ra  (hh e]rb  (hh"e]rc  (hhe]rd  (h%h&eeejR  jR  jR  jR  jR  jR  ]re  (h]rf  (h]rg  (h]rh  (hh	e]ri  (hh	e]rj  (hhe]rk  (h]rl  (hh	e]rm  (hhe]rn  (hhe]ro  (j�  ]rp  (hh	e]rq  (hheeee]rr  (hhee]rs  (h]rt  (hh e]ru  (hh"e]rv  (hhe]rw  (h%h&eeeje  je  ]rx  (h]ry  (h]rz  (h]r{  (hh	e]r|  (hh	e]r}  (hhe]r~  (h]r  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeejx  jx  jx  jx  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r 	  (hh	e]r	  (hh	e]r	  (hhe]r	  (h]r	  (hh	e]r	  (hhe]r	  (hhe]r	  (j�  ]r	  (hh	e]r		  (hheeee]r
	  (hhee]r	  (h]r	  (hh e]r	  (hh"e]r	  (hhe]r	  (h%h&eeej�  j�  j�  ]r	  (h]r	  (h]r	  (h]r	  (hh	e]r	  (hh	e]r	  (hhe]r	  (h]r	  (hh	e]r	  (hhe]r	  (hhe]r	  (j�  ]r	  (hh	e]r	  (hheeee]r	  (hhee]r	  (h]r	  (hh e]r 	  (hh"e]r!	  (hhe]r"	  (h%h&eeej	  ]r#	  (h]r$	  (h]r%	  (h]r&	  (hh	e]r'	  (hh	e]r(	  (hhe]r)	  (h]r*	  (hh	e]r+	  (hhe]r,	  (hhe]r-	  (j�  ]r.	  (hh	e]r/	  (hheeee]r0	  (hhee]r1	  (h]r2	  (hh e]r3	  (hh"e]r4	  (hhe]r5	  (h%h&eeej#	  j#	  j#	  ]r6	  (h]r7	  (h]r8	  (h]r9	  (hh	e]r:	  (hh	e]r;	  (hhe]r<	  (h]r=	  (hh	e]r>	  (hhe]r?	  (hhe]r@	  (j�  ]rA	  (hh	e]rB	  (hheeee]rC	  (hhee]rD	  (h]rE	  (hh e]rF	  (hh"e]rG	  (hhe]rH	  (h%h&eee]rI	  (h]rJ	  (h]rK	  (h]rL	  (hh	e]rM	  (hh	e]rN	  (hhe]rO	  (h]rP	  (hh	e]rQ	  (hhe]rR	  (hhe]rS	  (j�  ]rT	  (hh	e]rU	  (hheeee]rV	  (hhee]rW	  (h]rX	  (hh e]rY	  (hh"e]rZ	  (hhe]r[	  (h%h&eeejI	  jI	  ]r\	  (h]r]	  (h]r^	  (h]r_	  (hh	e]r`	  (hh	e]ra	  (hhe]rb	  (h]rc	  (hhe]rd	  (hhe]re	  (hhe]rf	  (j�  ]rg	  (hh	e]rh	  (hheeee]ri	  (hhee]rj	  (h]rk	  (hh e]rl	  (hh"e]rm	  (hhe]rn	  (h%h&eeej\	  j\	  j\	  j\	  j\	  j\	  j\	  j\	  j\	  ]ro	  (h]rp	  (h]rq	  (h]rr	  (hh	e]rs	  (hh	e]rt	  (hhe]ru	  (h]rv	  (hhe]rw	  (hhe]rx	  (hhe]ry	  (j�  ]rz	  (hh	e]r{	  (hheeee]r|	  (hhee]r}	  (h]r~	  (hh e]r	  (hh"e]r�	  (hhe]r�	  (h%h&eee]r�	  (h]r�	  (h]r�	  (h]r�	  (hh	e]r�	  (hh	e]r�	  (hhe]r�	  (h]r�	  (hhe]r�	  (hhe]r�	  (hhe]r�	  (j�  ]r�	  (hh	e]r�	  (hheeee]r�	  (hhee]r�	  (h]r�	  (hh e]r�	  (hh"e]r�	  (hhe]r�	  (h%h&eeej�	  j�	  j�	  j�	  j�	  ]r�	  (h]r�	  (h]r�	  (h]r�	  (hh	e]r�	  (hh	e]r�	  (hhe]r�	  (h]r�	  (hhe]r�	  (hhe]r�	  (hhe]r�	  (j�  ]r�	  (hh	e]r�	  (hheeee]r�	  (hhee]r�	  (h]r�	  (hh e]r�	  (hh"e]r�	  (hhe]r�	  (h%h&eeej�	  j�	  ]r�	  (h]r�	  (h]r�	  (h]r�	  (hh	e]r�	  (hh	e]r�	  (hhe]r�	  (h]r�	  (hhe]r�	  (hhe]r�	  (hhe]r�	  (j�  ]r�	  (hh	e]r�	  (hheeee]r�	  (hhee]r�	  (h]r�	  (hh e]r�	  (hh"e]r�	  (hhe]r�	  (h%h&eeej�	  j�	  j�	  ]r�	  (h]r�	  (h]r�	  (h]r�	  (hh	e]r�	  (hh	e]r�	  (hhe]r�	  (h]r�	  (hhe]r�	  (hhe]r�	  (hhe]r�	  (j�  ]r�	  (hh	e]r�	  (hheeee]r�	  (hhee]r�	  (h]r�	  (hh e]r�	  (hh"e]r�	  (hhe]r�	  (h%h&eeej�	  j�	  j�	  ]r�	  (h]r�	  (h]r�	  (h]r�	  (hh	e]r�	  (hh	e]r�	  (hhe]r�	  (h]r�	  (hhe]r�	  (hhe]r�	  (hhe]r�	  (j�  ]r�	  (hh	e]r�	  (hheeee]r�	  (hhee]r�	  (h]r�	  (hh e]r�	  (hh"e]r�	  (hhe]r�	  (h%h&eeej�	  j�	  j�	  ]r�	  (h]r�	  (h]r�	  (h]r�	  (hh	e]r�	  (hh	e]r�	  (hhe]r�	  (h]r�	  (hhe]r�	  (hhe]r�	  (hhe]r�	  (j�  ]r�	  (hh	e]r�	  (hheeee]r�	  (hhee]r�	  (h]r�	  (hh e]r�	  (hh"e]r�	  (hhe]r�	  (h%h&eeej�	  j�	  j�	  j�	  ]r�	  (h]r�	  (h]r�	  (h]r�	  (hh	e]r�	  (hh	e]r�	  (hhe]r�	  (h]r�	  (hhe]r�	  (hhe]r�	  (hhe]r�	  (j�  ]r�	  (hh	e]r 
  (hheeee]r
  (hhee]r
  (h]r
  (hh e]r
  (hh"e]r
  (hhe]r
  (h%h&eeej�	  j�	  ]r
  (h]r
  (h]r	
  (h]r

  (hh	e]r
  (hh	e]r
  (hhe]r
  (h]r
  (hhe]r
  (hhe]r
  (hhe]r
  (j�  ]r
  (hh	e]r
  (hheeee]r
  (hhee]r
  (h]r
  (hh e]r
  (hh"e]r
  (hhe]r
  (h%h&eeej
  j
  j
  ]r
  (h]r
  (h]r
  (h]r
  (hh	e]r
  (hh	e]r
  (hhe]r 
  (h]r!
  (hhe]r"
  (hhe]r#
  (hhe]r$
  (j�  ]r%
  (hh	e]r&
  (hheeee]r'
  (hhee]r(
  (h]r)
  (hh e]r*
  (hh"e]r+
  (hhe]r,
  (h%h&eee]r-
  (h]r.
  (h]r/
  (h]r0
  (hh	e]r1
  (hh	e]r2
  (hhe]r3
  (h]r4
  (hhe]r5
  (hhe]r6
  (hhe]r7
  (j�  ]r8
  (hh	e]r9
  (hheeee]r:
  (hhee]r;
  (h]r<
  (hh e]r=
  (hh"e]r>
  (hhe]r?
  (h%h&eee]r@
  (h]rA
  (h]rB
  (h]rC
  (hh	e]rD
  (hh	e]rE
  (hhe]rF
  (h]rG
  (hhe]rH
  (hhe]rI
  (hhe]rJ
  (j�  ]rK
  (hh	e]rL
  (hheeee]rM
  (hhee]rN
  (h]rO
  (hh e]rP
  (hh"e]rQ
  (hhe]rR
  (h%h&eeej@
  j@
  j@
  ]rS
  (h]rT
  (h]rU
  (h]rV
  (hh	e]rW
  (hh	e]rX
  (hhe]rY
  (h]rZ
  (hh	e]r[
  (hhe]r\
  (hhe]r]
  (j�  ]r^
  (hh	e]r_
  (hheeee]r`
  (hhee]ra
  (h]rb
  (hh e]rc
  (hh"e]rd
  (hhe]re
  (h%h&eee]rf
  (h]rg
  (h]rh
  (h]ri
  (hh	e]rj
  (hh	e]rk
  (hhe]rl
  (h]rm
  (hh	e]rn
  (hhe]ro
  (hhe]rp
  (j�  ]rq
  (hh	e]rr
  (hheeee]rs
  (hhee]rt
  (h]ru
  (hh e]rv
  (hh"e]rw
  (hhe]rx
  (h%h&eee]ry
  (h]rz
  (h]r{
  (h]r|
  (hh	e]r}
  (hh	e]r~
  (hhe]r
  (h]r�
  (hh	e]r�
  (hhe]r�
  (hhe]r�
  (j�  ]r�
  (hh	e]r�
  (hheeee]r�
  (hhee]r�
  (h]r�
  (hh e]r�
  (hh"e]r�
  (hhe]r�
  (h%h&eeejy
  jy
  jy
  jy
  jy
  jy
  jy
  ]r�
  (h]r�
  (h]r�
  (h]r�
  (hh	e]r�
  (hh	e]r�
  (hhe]r�
  (h]r�
  (hh	e]r�
  (hhe]r�
  (hhe]r�
  (j�  ]r�
  (hh	e]r�
  (hheeee]r�
  (hhee]r�
  (h]r�
  (hh e]r�
  (hh"e]r�
  (hhe]r�
  (h%h&eeej�
  j�
  j�
  j�
  j�
  ]r�
  (h]r�
  (h]r�
  (h]r�
  (hh	e]r�
  (hh	e]r�
  (hhe]r�
  (h]r�
  (hh	e]r�
  (hhe]r�
  (hhe]r�
  (j�  ]r�
  (hh	e]r�
  (hheeee]r�
  (hhee]r�
  (h]r�
  (hh e]r�
  (hh"e]r�
  (hhe]r�
  (h%h&eeej�
  j�
  j�
  ]r�
  (h]r�
  (h]r�
  (h]r�
  (hh	e]r�
  (hh	e]r�
  (hhe]r�
  (h]r�
  (hh	e]r�
  (hhe]r�
  (hhe]r�
  (j�  ]r�
  (hh	e]r�
  (hheeee]r�
  (hhee]r�
  (h]r�
  (hh e]r�
  (hh"e]r�
  (hhe]r�
  (h%h&eeej�
  j�
  j�
  ]r�
  (h]r�
  (h]r�
  (h]r�
  (hh	e]r�
  (hh	e]r�
  (hhe]r�
  (h]r�
  (hh	e]r�
  (hhe]r�
  (hhe]r�
  (j�  ]r�
  (hh	e]r�
  (hheeee]r�
  (hhee]r�
  (h]r�
  (hh e]r�
  (hh"e]r�
  (hhe]r�
  (h%h&eeej�
  j�
  j�
  j�
  j�
  j�
  ]r�
  (h]r�
  (h]r�
  (h]r�
  (hh	e]r�
  (hh	e]r�
  (hhe]r�
  (h]r�
  (hhe]r�
  (hhe]r�
  (hhe]r�
  (j�  ]r�
  (hh	e]r�
  (hheeee]r�
  (hhee]r�
  (h]r�
  (hh e]r�
  (hh"e]r�
  (hhe]r�
  (h%h&eee]r�
  (h]r�
  (h]r�
  (h]r�
  (hh	e]r�
  (hh	e]r�
  (hhe]r�
  (h]r�
  (hhe]r�
  (hhe]r�
  (hhe]r�
  (j�  ]r�
  (hh	e]r�
  (hheeee]r�
  (hhee]r�
  (h]r�
  (hh e]r�
  (hh"e]r�
  (hhe]r�
  (h%h&eeej�
  j�
  j�
  ]r�
  (h]r�
  (h]r   (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r  (hhe]r  (j�  ]r	  (hh	e]r
  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hhe]r  (h%h&eeej�
  j�
  j�
  j�
  j�
  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hh	e]r  (hhe]r  (hhe]r  (j�  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r   (hh e]r!  (hh"e]r"  (hhe]r#  (h%h&eee]r$  (h]r%  (h]r&  (h]r'  (hh	e]r(  (hh	e]r)  (hhe]r*  (h]r+  (hh	e]r,  (hhe]r-  (hhe]r.  (j�  ]r/  (hh	e]r0  (hheeee]r1  (hhee]r2  (h]r3  (hh e]r4  (hh"e]r5  (hhe]r6  (h%h&eeej$  j$  j$  j$  ]r7  (h]r8  (h]r9  (h]r:  (hh	e]r;  (hh	e]r<  (hhe]r=  (h]r>  (hh	e]r?  (hhe]r@  (hhe]rA  (j�  ]rB  (hh	e]rC  (hheeee]rD  (hhee]rE  (h]rF  (hh e]rG  (hh"e]rH  (hhe]rI  (h%h&eeej7  j7  j7  ]rJ  (h]rK  (h]rL  (h]rM  (hh	e]rN  (hh	e]rO  (hhe]rP  (h]rQ  (hh	e]rR  (hhe]rS  (hhe]rT  (j�  ]rU  (hh	e]rV  (hheeee]rW  (hhee]rX  (h]rY  (hh e]rZ  (hh"e]r[  (hhe]r\  (h%h&eee]r]  (h]r^  (h]r_  (h]r`  (hh	e]ra  (hh	e]rb  (hhe]rc  (h]rd  (hh	e]re  (hhe]rf  (hhe]rg  (j�  ]rh  (hh	e]ri  (hheeee]rj  (hhee]rk  (h]rl  (hh e]rm  (hh"e]rn  (hhe]ro  (h%h&eee]rp  (h]rq  (h]rr  (h]rs  (hh	e]rt  (hh	e]ru  (hhe]rv  (h]rw  (hh	e]rx  (hhe]ry  (hhe]rz  (j�  ]r{  (hh	e]r|  (hheeee]r}  (hhee]r~  (h]r  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeejp  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r   (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hhe]r  (h%h&eeej�  j�  j�  j�  j�  ]r  (h]r	  (h]r
  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hh	e]r  (hhe]r  (hhe]r  (j�  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hh	e]r  (h%h&eeej  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r   (hhe]r!  (h]r"  (hh	e]r#  (hhe]r$  (hhe]r%  (j�  ]r&  (hh	e]r'  (hheeee]r(  (hhee]r)  (h]r*  (hh e]r+  (hh"e]r,  (hh	e]r-  (h%h&eeej  ]r.  (h]r/  (h]r0  (h]r1  (hh	e]r2  (hh	e]r3  (hhe]r4  (h]r5  (hh	e]r6  (hhe]r7  (hhe]r8  (j�  ]r9  (hh	e]r:  (hheeee]r;  (hhee]r<  (h]r=  (hh e]r>  (hh"e]r?  (hhe]r@  (h%h&eeej.  j.  j.  j.  j.  j.  ]rA  (h]rB  (h]rC  (h]rD  (hh	e]rE  (hh	e]rF  (hhe]rG  (h]rH  (hh	e]rI  (hhe]rJ  (hhe]rK  (j�  ]rL  (hh	e]rM  (hheeee]rN  (hhee]rO  (h]rP  (hh e]rQ  (hh"e]rR  (hhe]rS  (h%h&eeejA  ]rT  (h]rU  (h]rV  (h]rW  (hh	e]rX  (hh	e]rY  (hhe]rZ  (h]r[  (hhe]r\  (hhe]r]  (hhe]r^  (j�  ]r_  (hh	e]r`  (hheeee]ra  (hhee]rb  (h]rc  (hh e]rd  (hh"e]re  (hhe]rf  (h%h&eeejT  jT  ]rg  (h]rh  (h]ri  (h]rj  (hh	e]rk  (hh	e]rl  (hhe]rm  (h]rn  (hhe]ro  (hhe]rp  (hhe]rq  (j�  ]rr  (hh	e]rs  (hheeee]rt  (hhee]ru  (h]rv  (hh e]rw  (hh"e]rx  (hhe]ry  (h%h&eeejg  ]rz  (h]r{  (h]r|  (h]r}  (hh	e]r~  (hh	e]r  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeejz  jz  jz  jz  jz  jz  jz  jz  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  ]r�  (h]r   (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r  (hhe]r	  (j�  ]r
  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hh	e]r  (h%h&eeej�  j�  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r  (hhe]r  (j�  ]r  (hh	e]r  (hheeee]r  (hhee]r   (h]r!  (hh e]r"  (hh"e]r#  (hh	e]r$  (h%h&eeej  j  j  ]r%  (h]r&  (h]r'  (h]r(  (hh	e]r)  (hh	e]r*  (hhe]r+  (h]r,  (hh	e]r-  (hhe]r.  (hhe]r/  (j�  ]r0  (hh	e]r1  (hheeee]r2  (hhee]r3  (h]r4  (hh e]r5  (hh"e]r6  (hh	e]r7  (h%h&eee]r8  (h]r9  (h]r:  (h]r;  (hh	e]r<  (hh	e]r=  (hhe]r>  (h]r?  (hh	e]r@  (hhe]rA  (hhe]rB  (j�  ]rC  (hh	e]rD  (hheeee]rE  (hhee]rF  (h]rG  (hh e]rH  (hh"e]rI  (hh	e]rJ  (h%h&eeej8  j8  j8  j8  j8  j8  j8  j8  j8  j8  j8  j8  ]rK  (h]rL  (h]rM  (h]rN  (hh	e]rO  (hh	e]rP  (hhe]rQ  (h]rR  (hh	e]rS  (hhe]rT  (hhe]rU  (j�  ]rV  (hh	e]rW  (hheeee]rX  (hhee]rY  (h]rZ  (hh e]r[  (hh"e]r\  (hh	e]r]  (h%h&eeejK  jK  jK  jK  jK  jK  jK  ]r^  (h]r_  (h]r`  (h]ra  (hh	e]rb  (hh	e]rc  (hhe]rd  (h]re  (hh	e]rf  (hhe]rg  (hhe]rh  (j�  ]ri  (hh	e]rj  (hheeee]rk  (hhee]rl  (h]rm  (hh e]rn  (hh"e]ro  (hh	e]rp  (h%h&eeej^  j^  ]rq  (h]rr  (h]rs  (h]rt  (hh	e]ru  (hh	e]rv  (hhe]rw  (h]rx  (hh	e]ry  (hhe]rz  (hhe]r{  (j�  ]r|  (hh	e]r}  (hheeee]r~  (hhee]r  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeejq  jq  jq  jq  jq  jq  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r   (X	   Next-Mover  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hh	e]r	  (h%h&eee]r
  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r  (hhe]r  (j  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hh	e]r  (h%h&eeej
  ]r  (h]r  (h]r  (h]r   (hh	e]r!  (hh	e]r"  (hhe]r#  (h]r$  (hhe]r%  (hhe]r&  (hhe]r'  (j  ]r(  (hh	e]r)  (hheeee]r*  (hhee]r+  (h]r,  (hh e]r-  (hh"e]r.  (hh	e]r/  (h%h&eeej  ]r0  (h]r1  (h]r2  (h]r3  (hh	e]r4  (hh	e]r5  (hhe]r6  (h]r7  (hhe]r8  (hhe]r9  (hhe]r:  (j  ]r;  (hh	e]r<  (hheeee]r=  (hhee]r>  (h]r?  (hh e]r@  (hh"e]rA  (hh	e]rB  (h%h&eee]rC  (h]rD  (h]rE  (h]rF  (hh	e]rG  (hh	e]rH  (hhe]rI  (h]rJ  (hhe]rK  (hhe]rL  (hhe]rM  (j  ]rN  (hh	e]rO  (hheeee]rP  (hhee]rQ  (h]rR  (hh e]rS  (hh"e]rT  (hh	e]rU  (h%h&eeejC  jC  jC  jC  jC  jC  jC  jC  jC  jC  jC  jC  jC  jC  ]rV  (h]rW  (h]rX  (h]rY  (hh	e]rZ  (hh	e]r[  (hhe]r\  (h]r]  (hhe]r^  (hhe]r_  (hhe]r`  (j  ]ra  (hh	e]rb  (hheeee]rc  (hhee]rd  (h]re  (hh e]rf  (hh"e]rg  (hh	e]rh  (h%h&eee]ri  (h]rj  (h]rk  (h]rl  (hh	e]rm  (hh	e]rn  (hhe]ro  (h]rp  (hhe]rq  (hhe]rr  (hhe]rs  (j  ]rt  (hh	e]ru  (hheeee]rv  (hhee]rw  (h]rx  (hh e]ry  (hh"e]rz  (hh	e]r{  (h%h&eeeji  ji  ]r|  (h]r}  (h]r~  (h]r  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r   (h%h&eeej�  j�  j�  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hhe]r	  (hhe]r
  (hhe]r  (j  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hh	e]r  (h%h&eeej  j  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r  (hhe]r  (j  ]r  (hh	e]r   (hheeee]r!  (hhee]r"  (h]r#  (hh e]r$  (hh"e]r%  (hh	e]r&  (h%h&eeej  j  j  j  j  j  j  ]r'  (h]r(  (h]r)  (h]r*  (hh	e]r+  (hh	e]r,  (hhe]r-  (h]r.  (hhe]r/  (hhe]r0  (hhe]r1  (j  ]r2  (hh	e]r3  (hheeee]r4  (hhee]r5  (h]r6  (hh e]r7  (hh"e]r8  (hh	e]r9  (h%h&eeej'  ]r:  (h]r;  (h]r<  (h]r=  (hh	e]r>  (hh	e]r?  (hhe]r@  (h]rA  (hhe]rB  (hhe]rC  (hhe]rD  (j  ]rE  (hh	e]rF  (hheeee]rG  (hhee]rH  (h]rI  (hh e]rJ  (hh"e]rK  (hh	e]rL  (h%h&eeej:  j:  j:  ]rM  (h]rN  (h]rO  (h]rP  (hh	e]rQ  (hh	e]rR  (hhe]rS  (h]rT  (hhe]rU  (hhe]rV  (hhe]rW  (j  ]rX  (hh	e]rY  (hheeee]rZ  (hhee]r[  (h]r\  (hh e]r]  (hh"e]r^  (hh	e]r_  (h%h&eeejM  jM  ]r`  (h]ra  (h]rb  (h]rc  (hh	e]rd  (hh	e]re  (hhe]rf  (h]rg  (hhe]rh  (hhe]ri  (hhe]rj  (j  ]rk  (hh	e]rl  (hheeee]rm  (hhee]rn  (h]ro  (hh e]rp  (hh"e]rq  (hh	e]rr  (h%h&eee]rs  (h]rt  (h]ru  (h]rv  (hh	e]rw  (hh	e]rx  (hhe]ry  (h]rz  (hhe]r{  (hhe]r|  (hhe]r}  (j  ]r~  (hh	e]r  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeejs  js  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r   (hhe]r  (hhe]r  (j  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r	  (hh	e]r
  (h%h&eeej�  j�  j�  j�  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r  (hhe]r  (j  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hh	e]r  (h%h&eee]r  (h]r  (h]r   (h]r!  (hh	e]r"  (hh	e]r#  (hhe]r$  (h]r%  (hhe]r&  (hhe]r'  (hhe]r(  (j  ]r)  (hh	e]r*  (hheeee]r+  (hhee]r,  (h]r-  (hh e]r.  (hh"e]r/  (hh	e]r0  (h%h&eeej  j  j  ]r1  (h]r2  (h]r3  (h]r4  (hh	e]r5  (hh	e]r6  (hhe]r7  (h]r8  (hhe]r9  (hhe]r:  (hhe]r;  (j  ]r<  (hh	e]r=  (hheeee]r>  (hhee]r?  (h]r@  (hh e]rA  (hh"e]rB  (hh	e]rC  (h%h&eeej1  j1  ]rD  (h]rE  (h]rF  (h]rG  (hh	e]rH  (hh	e]rI  (hhe]rJ  (h]rK  (hhe]rL  (hhe]rM  (hhe]rN  (j  ]rO  (hh	e]rP  (hheeee]rQ  (hhee]rR  (h]rS  (hh e]rT  (hh"e]rU  (hh	e]rV  (h%h&eeejD  jD  jD  jD  ]rW  (h]rX  (h]rY  (h]rZ  (hh	e]r[  (hh	e]r\  (hhe]r]  (h]r^  (hhe]r_  (hhe]r`  (hhe]ra  (j  ]rb  (hh	e]rc  (hheeee]rd  (hhee]re  (h]rf  (hh e]rg  (hh"e]rh  (hh	e]ri  (h%h&eeejW  jW  jW  jW  ]rj  (h]rk  (h]rl  (h]rm  (hh	e]rn  (hh	e]ro  (hhe]rp  (h]rq  (hhe]rr  (hhe]rs  (hhe]rt  (j  ]ru  (hh	e]rv  (hheeee]rw  (hhee]rx  (h]ry  (hh e]rz  (hh"e]r{  (hh	e]r|  (h%h&eeejj  ]r}  (h]r~  (h]r  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej}  j}  j}  j}  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hh	e]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r   (hhe]r  (h%h&eeej�  j�  j�  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r	  (hhe]r
  (hhe]r  (hhe]r  (j  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hh	e]r  (h%h&eeej  j  j  j  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hhe]r  (hhe]r  (hhe]r  (j  ]r   (hh	e]r!  (hheeee]r"  (hhee]r#  (h]r$  (hh e]r%  (hh"e]r&  (hh	e]r'  (h%h&eeej  j  j  ]r(  (h]r)  (h]r*  (h]r+  (hh	e]r,  (hh	e]r-  (hhe]r.  (h]r/  (hhe]r0  (hhe]r1  (hhe]r2  (j  ]r3  (hh	e]r4  (hheeee]r5  (hhee]r6  (h]r7  (hh e]r8  (hh"e]r9  (hh	e]r:  (h%h&eeej(  j(  ]r;  (h]r<  (h]r=  (h]r>  (hh	e]r?  (hh	e]r@  (hhe]rA  (h]rB  (hhe]rC  (hhe]rD  (hhe]rE  (j  ]rF  (hh	e]rG  (hheeee]rH  (hhee]rI  (h]rJ  (hh e]rK  (hh"e]rL  (hh	e]rM  (h%h&eeej;  j;  j;  ]rN  (h]rO  (h]rP  (h]rQ  (hh	e]rR  (hh	e]rS  (hhe]rT  (h]rU  (hhe]rV  (hhe]rW  (hhe]rX  (j  ]rY  (hh	e]rZ  (hheeee]r[  (hhee]r\  (h]r]  (hh e]r^  (hh"e]r_  (hhe]r`  (h%h&eeejN  jN  jN  ]ra  (h]rb  (h]rc  (h]rd  (hh	e]re  (hh	e]rf  (hhe]rg  (h]rh  (hhe]ri  (hhe]rj  (hhe]rk  (j  ]rl  (hh	e]rm  (hheeee]rn  (hhee]ro  (h]rp  (hh e]rq  (hh"e]rr  (hhe]rs  (h%h&eeeja  ja  ja  ]rt  (h]ru  (h]rv  (h]rw  (hh	e]rx  (hh	e]ry  (hhe]rz  (h]r{  (hhe]r|  (hhe]r}  (hhe]r~  (j  ]r  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeejt  jt  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eee]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hhe]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r�  (hh	e]r�  (hhe]r�  (hhe]r�  (j  ]r�  (hh	e]r�  (hheeee]r�  (hhee]r�  (h]r�  (hh e]r�  (hh"e]r�  (hhe]r�  (h%h&eeej�  ]r�  (h]r�  (h]r�  (h]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (h]r   (hh	e]r  (hhe]r  (hhe]r  (j  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r	  (hh"e]r
  (hhe]r  (h%h&eeej�  j�  ]r  (h]r  (h]r  (h]r  (hh	e]r  (hh	e]r  (hhe]r  (h]r  (hh	e]r  (hhe]r  (hhe]r  (j  ]r  (hh	e]r  (hheeee]r  (hhee]r  (h]r  (hh e]r  (hh"e]r  (hhe]r  (h%h&eeej  j  j  j  j  j  j  j  j  ]r  (h]r   (h]r!  (h]r"  (hh	e]r#  (hh	e]r$  (hhe]r%  (h]r&  (hh	e]r'  (hhe]r(  (hhe]r)  (j  ]r*  (hh	e]r+  (hheeee]r,  (hhee]r-  (h]r.  (hh e]r/  (hh"e]r0  (hhe]r1  (h%h&eee]r2  (h]r3  (h]r4  (h]r5  (hh	e]r6  (hh	e]r7  (hhe]r8  (h]r9  (hhe]r:  (hhe]r;  (hhe]r<  (j  ]r=  (hh	e]r>  (hheeee]r?  (hhee]r@  (h]rA  (hh e]rB  (hh"e]rC  (hhe]rD  (h%h&eeee(]rE  (X   NormrF  ]rG  (X   OblrH  ]rI  (X   MovedrJ  ]rK  (hh	e]rL  (hhe]rM  (hX   1rN  e]rO  (X   MovedrP  ]rQ  (hh	e]rR  (hh	e]rS  (hhe]rT  (X	   Next-MoverU  ]rV  (hhe]rW  (hheeee]rX  (hheee]rY  (jF  ]rZ  (jH  ]r[  (jJ  ]r\  (hh	e]r]  (hhe]r^  (hjN  e]r_  (jP  ]r`  (hh	e]ra  (hh	e]rb  (hhe]rc  (jU  ]rd  (hhe]re  (hheeee]rf  (hheeejY  jY  jY  jY  jY  jY  jY  jY  jY  jY  jY  jY  jY  jY  jY  ]rg  (jF  ]rh  (jH  ]ri  (jJ  ]rj  (hh	e]rk  (hhe]rl  (hjN  e]rm  (jP  ]rn  (hh	e]ro  (hh	e]rp  (hhe]rq  (jU  ]rr  (hhe]rs  (hheeee]rt  (hheee]ru  (jF  ]rv  (jH  ]rw  (jJ  ]rx  (hh	e]ry  (hhe]rz  (hjN  e]r{  (jP  ]r|  (hh	e]r}  (hh	e]r~  (hhe]r  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r   (hheeej�  j�  j�  j�  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (jP  ]r  (hh	e]r	  (hh	e]r
  (hhe]r  (jU  ]r  (hhe]r  (hheeee]r  (hheeej  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (jP  ]r  (hh	e]r  (hh	e]r  (hhe]r  (jU  ]r  (hhe]r  (hheeee]r  (hheeej  ]r  (jF  ]r  (jH  ]r  (jJ  ]r   (hh"e]r!  (hhe]r"  (hjN  e]r#  (jP  ]r$  (hh	e]r%  (hh	e]r&  (hhe]r'  (jU  ]r(  (hhe]r)  (hheeee]r*  (hheeej  j  ]r+  (jF  ]r,  (jH  ]r-  (jJ  ]r.  (hh"e]r/  (hhe]r0  (hjN  e]r1  (jP  ]r2  (hh	e]r3  (hh	e]r4  (hhe]r5  (jU  ]r6  (hhe]r7  (hheeee]r8  (hheee]r9  (jF  ]r:  (jH  ]r;  (jJ  ]r<  (hh"e]r=  (hhe]r>  (hjN  e]r?  (jP  ]r@  (hh	e]rA  (hh	e]rB  (hhe]rC  (jU  ]rD  (hhe]rE  (hheeee]rF  (hheee]rG  (jF  ]rH  (jH  ]rI  (jJ  ]rJ  (hh"e]rK  (hhe]rL  (hjN  e]rM  (jP  ]rN  (hh	e]rO  (hh	e]rP  (hhe]rQ  (jU  ]rR  (hhe]rS  (hheeee]rT  (hheeejG  jG  jG  jG  ]rU  (jF  ]rV  (jH  ]rW  (jJ  ]rX  (hh"e]rY  (hh	e]rZ  (hjN  e]r[  (jP  ]r\  (hh	e]r]  (hh	e]r^  (hhe]r_  (jU  ]r`  (hhe]ra  (hheeee]rb  (hheeejU  jU  jU  ]rc  (jF  ]rd  (jH  ]re  (jJ  ]rf  (hh"e]rg  (hh	e]rh  (hjN  e]ri  (jP  ]rj  (hh	e]rk  (hh	e]rl  (hhe]rm  (jU  ]rn  (hhe]ro  (hheeee]rp  (hheeejc  jc  jc  jc  jc  jc  ]rq  (jF  ]rr  (jH  ]rs  (jJ  ]rt  (hh"e]ru  (hh	e]rv  (hjN  e]rw  (jP  ]rx  (hh	e]ry  (hh	e]rz  (hhe]r{  (jU  ]r|  (hhe]r}  (hheeee]r~  (hheeejq  jq  jq  ]r  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hh	e]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej  j  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hh	e]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hh	e]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hh	e]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hh	e]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hh	e]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hh	e]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hh	e]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hh	e]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r   (hh"e]r  (hhe]r  (hjN  e]r  (jP  ]r  (hh	e]r  (hh	e]r  (hhe]r  (jU  ]r  (hhe]r	  (hheeee]r
  (hheeej�  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (jP  ]r  (hh	e]r  (hh	e]r  (hhe]r  (jU  ]r  (hhe]r  (hheeee]r  (hheee]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (jP  ]r   (hh	e]r!  (hh	e]r"  (hhe]r#  (jU  ]r$  (hhe]r%  (hheeee]r&  (hheee]r'  (jF  ]r(  (jH  ]r)  (jJ  ]r*  (hh"e]r+  (hhe]r,  (hjN  e]r-  (jP  ]r.  (hh	e]r/  (hh	e]r0  (hhe]r1  (jU  ]r2  (hhe]r3  (hheeee]r4  (hheeej'  j'  j'  ]r5  (jF  ]r6  (jH  ]r7  (jJ  ]r8  (hh"e]r9  (hhe]r:  (hjN  e]r;  (jP  ]r<  (hh	e]r=  (hh	e]r>  (hhe]r?  (jU  ]r@  (hhe]rA  (hheeee]rB  (hheeej5  j5  j5  j5  j5  j5  j5  j5  j5  j5  j5  j5  ]rC  (jF  ]rD  (jH  ]rE  (jJ  ]rF  (hh"e]rG  (hhe]rH  (hjN  e]rI  (jP  ]rJ  (hh	e]rK  (hh	e]rL  (hhe]rM  (jU  ]rN  (hhe]rO  (hheeee]rP  (hheee]rQ  (jF  ]rR  (jH  ]rS  (jJ  ]rT  (hh"e]rU  (hhe]rV  (hjN  e]rW  (jP  ]rX  (hh	e]rY  (hh	e]rZ  (hhe]r[  (jU  ]r\  (hhe]r]  (hheeee]r^  (hheeejQ  ]r_  (jF  ]r`  (jH  ]ra  (jJ  ]rb  (hh"e]rc  (hhe]rd  (hjN  e]re  (jP  ]rf  (hh	e]rg  (hh	e]rh  (hhe]ri  (jU  ]rj  (hhe]rk  (hheeee]rl  (hheeej_  j_  j_  ]rm  (jF  ]rn  (jH  ]ro  (jJ  ]rp  (hh"e]rq  (hhe]rr  (hjN  e]rs  (jP  ]rt  (hh	e]ru  (hh	e]rv  (hhe]rw  (jU  ]rx  (hhe]ry  (hheeee]rz  (hheee]r{  (jF  ]r|  (jH  ]r}  (jJ  ]r~  (hh"e]r  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej{  j{  j{  j{  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r   (hh	e]r  (hh	e]r  (hhe]r  (jU  ]r  (hhe]r  (hheeee]r  (hheeej�  j�  ]r  (jF  ]r  (jH  ]r	  (jJ  ]r
  (hh"e]r  (hhe]r  (hjN  e]r  (jP  ]r  (hh	e]r  (hh	e]r  (hhe]r  (jU  ]r  (hhe]r  (hheeee]r  (hheee]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (jP  ]r  (hh	e]r  (hh	e]r  (hhe]r  (jU  ]r   (hhe]r!  (hheeee]r"  (hheeej  ]r#  (jF  ]r$  (jH  ]r%  (jJ  ]r&  (hh"e]r'  (hhe]r(  (hjN  e]r)  (jP  ]r*  (hh	e]r+  (hh	e]r,  (hhe]r-  (jU  ]r.  (hhe]r/  (hheeee]r0  (hheeej#  j#  j#  j#  j#  ]r1  (jF  ]r2  (jH  ]r3  (jJ  ]r4  (hh"e]r5  (hhe]r6  (hjN  e]r7  (jP  ]r8  (hh	e]r9  (hh	e]r:  (hhe]r;  (jU  ]r<  (hhe]r=  (hheeee]r>  (hheeej1  ]r?  (jF  ]r@  (jH  ]rA  (jJ  ]rB  (hh"e]rC  (hhe]rD  (hjN  e]rE  (jP  ]rF  (hh	e]rG  (hh	e]rH  (hhe]rI  (jU  ]rJ  (hhe]rK  (hheeee]rL  (hheeej?  j?  j?  j?  ]rM  (jF  ]rN  (jH  ]rO  (jJ  ]rP  (hh"e]rQ  (hhe]rR  (hjN  e]rS  (jP  ]rT  (hh	e]rU  (hh	e]rV  (hhe]rW  (jU  ]rX  (hhe]rY  (hheeee]rZ  (hheeejM  jM  jM  ]r[  (jF  ]r\  (jH  ]r]  (jJ  ]r^  (hh"e]r_  (hhe]r`  (hjN  e]ra  (jP  ]rb  (hh	e]rc  (hh	e]rd  (hhe]re  (jU  ]rf  (hhe]rg  (hheeee]rh  (hheeej[  ]ri  (jF  ]rj  (jH  ]rk  (jJ  ]rl  (hh"e]rm  (hhe]rn  (hjN  e]ro  (jP  ]rp  (hh	e]rq  (hh	e]rr  (hhe]rs  (jU  ]rt  (hhe]ru  (hheeee]rv  (hheeeji  ji  ]rw  (jF  ]rx  (jH  ]ry  (jJ  ]rz  (hh"e]r{  (hhe]r|  (hjN  e]r}  (jP  ]r~  (hh	e]r  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeejw  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r�  (hhe]r�  (hheeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (jP  ]r�  (hh	e]r�  (hh	e]r�  (hhe]r�  (jU  ]r   (hhe]r  (hheeee]r  (hheee]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r  (hhe]r  (hjN  e]r	  (jP  ]r
  (hh	e]r  (hh	e]r  (hhe]r  (jU  ]r  (hhe]r  (hheeee]r  (hheeej  j  j  j  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r  (hh	e]r  (hjN  e]r  (jP  ]r  (hh	e]r  (hh	e]r  (hhe]r  (jU  ]r  (hhe]r  (hheeee]r  (hheeej  ]r  (jF  ]r   (jH  ]r!  (jJ  ]r"  (hh"e]r#  (hh	e]r$  (hjN  e]r%  (jP  ]r&  (hh	e]r'  (hh	e]r(  (hhe]r)  (jU  ]r*  (hhe]r+  (hheeee]r,  (hheeej  ]r-  (jF  ]r.  (jH  ]r/  (jJ  ]r0  (hh"e]r1  (hh	e]r2  (hjN  e]r3  (jP  ]r4  (hh	e]r5  (hh	e]r6  (hhe]r7  (jU  ]r8  (hhe]r9  (hheeee]r:  (hheeej-  j-  j-  j-  j-  j-  j-  j-  ]r;  (jF  ]r<  (jH  ]r=  (jJ  ]r>  (hh"e]r?  (hh	e]r@  (hjN  e]rA  (jP  ]rB  (hh	e]rC  (hh	e]rD  (hhe]rE  (jU  ]rF  (hhe]rG  (hheeee]rH  (hheeej;  j;  j;  j;  j;  j;  j;  j;  ]rI  (jF  ]rJ  (jH  ]rK  (jJ  ]rL  (hh"e]rM  (hh	e]rN  (hjN  e]rO  (jP  ]rP  (hh	e]rQ  (hh	e]rR  (hhe]rS  (jU  ]rT  (hhe]rU  (hheeee]rV  (hheeejI  jI  jI  jI  ]rW  (jF  ]rX  (jH  ]rY  (jJ  ]rZ  (hh"e]r[  (hh	e]r\  (hjN  e]r]  (X   Movedr^  ]r_  (hhe]r`  (hh	e]ra  (hhe]rb  (X	   Next-Moverc  ]rd  (hh	e]re  (hh	eeee]rf  (hheeejW  jW  jW  jW  jW  jW  jW  jW  ]rg  (jF  ]rh  (jH  ]ri  (jJ  ]rj  (hh"e]rk  (hhe]rl  (hjN  e]rm  (j^  ]rn  (hhe]ro  (hh	e]rp  (hhe]rq  (jc  ]rr  (hh	e]rs  (hh	eeee]rt  (hheeejg  jg  jg  jg  ]ru  (jF  ]rv  (jH  ]rw  (jJ  ]rx  (hh"e]ry  (hhe]rz  (hjN  e]r{  (j^  ]r|  (hhe]r}  (hh	e]r~  (hhe]r  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeeju  ju  ju  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r   (hheeej�  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh	e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r	  (hh	e]r
  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheee]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh	e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheeej  j  j  j  j  j  j  j  ]r  (jF  ]r  (jH  ]r  (jJ  ]r   (hh	e]r!  (hhe]r"  (hjN  e]r#  (j^  ]r$  (hhe]r%  (hh	e]r&  (hhe]r'  (jc  ]r(  (hh	e]r)  (hh	eeee]r*  (hheeej  j  j  j  j  ]r+  (jF  ]r,  (jH  ]r-  (jJ  ]r.  (hh	e]r/  (hhe]r0  (hjN  e]r1  (j^  ]r2  (hhe]r3  (hh	e]r4  (hhe]r5  (jc  ]r6  (hh	e]r7  (hh	eeee]r8  (hheeej+  j+  ]r9  (jF  ]r:  (jH  ]r;  (jJ  ]r<  (hh"e]r=  (hhe]r>  (hjN  e]r?  (j^  ]r@  (hhe]rA  (hh	e]rB  (hhe]rC  (jc  ]rD  (hh	e]rE  (hh	eeee]rF  (hheeej9  j9  j9  j9  ]rG  (jF  ]rH  (jH  ]rI  (jJ  ]rJ  (hh"e]rK  (hhe]rL  (hjN  e]rM  (j^  ]rN  (hhe]rO  (hh	e]rP  (hhe]rQ  (jc  ]rR  (hh	e]rS  (hh	eeee]rT  (hheeejG  jG  ]rU  (jF  ]rV  (jH  ]rW  (jJ  ]rX  (hh"e]rY  (hhe]rZ  (hjN  e]r[  (j^  ]r\  (hhe]r]  (hh	e]r^  (hhe]r_  (jc  ]r`  (hh	e]ra  (hh	eeee]rb  (hheee]rc  (jF  ]rd  (jH  ]re  (jJ  ]rf  (hh"e]rg  (hhe]rh  (hjN  e]ri  (j^  ]rj  (hhe]rk  (hh	e]rl  (hhe]rm  (jc  ]rn  (hh	e]ro  (hh	eeee]rp  (hheee]rq  (jF  ]rr  (jH  ]rs  (jJ  ]rt  (hh"e]ru  (hhe]rv  (hjN  e]rw  (j^  ]rx  (hhe]ry  (hh	e]rz  (hhe]r{  (jc  ]r|  (hh	e]r}  (hh	eeee]r~  (hheee]r  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r   (hh	e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r	  (hh	eeee]r
  (hheee]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh	e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheee]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh	e]r  (hhe]r  (hjN  e]r  (j^  ]r   (hhe]r!  (hh	e]r"  (hhe]r#  (jc  ]r$  (hh	e]r%  (hh	eeee]r&  (hheeej  j  j  j  j  j  j  j  j  j  j  ]r'  (jF  ]r(  (jH  ]r)  (jJ  ]r*  (hh"e]r+  (hhe]r,  (hjN  e]r-  (j^  ]r.  (hhe]r/  (hh	e]r0  (hhe]r1  (jc  ]r2  (hh	e]r3  (hh	eeee]r4  (hheeej'  j'  j'  j'  j'  ]r5  (jF  ]r6  (jH  ]r7  (jJ  ]r8  (hh	e]r9  (hhe]r:  (hjN  e]r;  (j^  ]r<  (hhe]r=  (hh	e]r>  (hhe]r?  (jc  ]r@  (hh	e]rA  (hh	eeee]rB  (hheeej5  j5  j5  ]rC  (jF  ]rD  (jH  ]rE  (jJ  ]rF  (hh	e]rG  (hhe]rH  (hjN  e]rI  (j^  ]rJ  (hhe]rK  (hh	e]rL  (hhe]rM  (jc  ]rN  (hh	e]rO  (hh	eeee]rP  (hheeejC  ]rQ  (jF  ]rR  (jH  ]rS  (jJ  ]rT  (hh	e]rU  (hhe]rV  (hjN  e]rW  (j^  ]rX  (hhe]rY  (hh	e]rZ  (hhe]r[  (jc  ]r\  (hh	e]r]  (hh	eeee]r^  (hheeejQ  jQ  jQ  jQ  jQ  jQ  ]r_  (jF  ]r`  (jH  ]ra  (jJ  ]rb  (hh	e]rc  (hhe]rd  (hjN  e]re  (j^  ]rf  (hhe]rg  (hh	e]rh  (hhe]ri  (jc  ]rj  (hh	e]rk  (hh	eeee]rl  (hheeej_  ]rm  (jF  ]rn  (jH  ]ro  (jJ  ]rp  (hh	e]rq  (hhe]rr  (hjN  e]rs  (j^  ]rt  (hhe]ru  (hh	e]rv  (hhe]rw  (jc  ]rx  (hh	e]ry  (hh	eeee]rz  (hheeejm  jm  jm  jm  jm  jm  jm  jm  jm  jm  jm  jm  jm  jm  jm  jm  ]r{  (jF  ]r|  (jH  ]r}  (jJ  ]r~  (hh	e]r  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r   (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheeej�  j�  ]r  (jF  ]r  (jH  ]r	  (jJ  ]r
  (hh	e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheeej  j  j  j  j  j  j  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh	e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r   (hh	e]r!  (hh	eeee]r"  (hheeej  j  j  j  ]r#  (jF  ]r$  (jH  ]r%  (jJ  ]r&  (hh"e]r'  (hhe]r(  (hjN  e]r)  (j^  ]r*  (hhe]r+  (hh	e]r,  (hhe]r-  (jc  ]r.  (hh	e]r/  (hh	eeee]r0  (hheeej#  j#  j#  j#  ]r1  (jF  ]r2  (jH  ]r3  (jJ  ]r4  (hh"e]r5  (hhe]r6  (hjN  e]r7  (j^  ]r8  (hhe]r9  (hh	e]r:  (hhe]r;  (jc  ]r<  (hh	e]r=  (hh	eeee]r>  (hheeej1  j1  ]r?  (jF  ]r@  (jH  ]rA  (jJ  ]rB  (hh	e]rC  (hhe]rD  (hjN  e]rE  (j^  ]rF  (hhe]rG  (hh	e]rH  (hhe]rI  (jc  ]rJ  (hh	e]rK  (hh	eeee]rL  (hheeej?  j?  ]rM  (jF  ]rN  (jH  ]rO  (jJ  ]rP  (hh	e]rQ  (hhe]rR  (hjN  e]rS  (j^  ]rT  (hhe]rU  (hh	e]rV  (hhe]rW  (jc  ]rX  (hh	e]rY  (hh	eeee]rZ  (hheeejM  ]r[  (jF  ]r\  (jH  ]r]  (jJ  ]r^  (hh"e]r_  (hhe]r`  (hjN  e]ra  (j^  ]rb  (hhe]rc  (hh	e]rd  (hhe]re  (jc  ]rf  (hh	e]rg  (hh	eeee]rh  (hheeej[  j[  ]ri  (jF  ]rj  (jH  ]rk  (jJ  ]rl  (hh"e]rm  (hhe]rn  (hjN  e]ro  (j^  ]rp  (hhe]rq  (hh	e]rr  (hhe]rs  (jc  ]rt  (hh	e]ru  (hh	eeee]rv  (hheeeji  ji  ]rw  (jF  ]rx  (jH  ]ry  (jJ  ]rz  (hh"e]r{  (hhe]r|  (hjN  e]r}  (j^  ]r~  (hhe]r  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeejw  jw  jw  jw  jw  jw  jw  jw  jw  jw  jw  jw  jw  jw  jw  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r   (hh	e]r  (hh	eeee]r  (hheee]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh	e]r  (hhe]r  (hjN  e]r	  (j^  ]r
  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheee]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh	e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheeej  ]r  (jF  ]r   (jH  ]r!  (jJ  ]r"  (hh	e]r#  (hhe]r$  (hjN  e]r%  (j^  ]r&  (hhe]r'  (hh	e]r(  (hhe]r)  (jc  ]r*  (hh	e]r+  (hh	eeee]r,  (hheeej  j  j  j  ]r-  (jF  ]r.  (jH  ]r/  (jJ  ]r0  (hh	e]r1  (hhe]r2  (hjN  e]r3  (j^  ]r4  (hhe]r5  (hh	e]r6  (hhe]r7  (jc  ]r8  (hh	e]r9  (hh	eeee]r:  (hheeej-  j-  j-  ]r;  (jF  ]r<  (jH  ]r=  (jJ  ]r>  (hh	e]r?  (hhe]r@  (hjN  e]rA  (j^  ]rB  (hhe]rC  (hh	e]rD  (hhe]rE  (jc  ]rF  (hh	e]rG  (hh	eeee]rH  (hheeej;  j;  j;  j;  ]rI  (jF  ]rJ  (jH  ]rK  (jJ  ]rL  (hh	e]rM  (hhe]rN  (hjN  e]rO  (j^  ]rP  (hhe]rQ  (hh	e]rR  (hhe]rS  (jc  ]rT  (hh	e]rU  (hh	eeee]rV  (hheeejI  jI  jI  ]rW  (jF  ]rX  (jH  ]rY  (jJ  ]rZ  (hh	e]r[  (hhe]r\  (hjN  e]r]  (j^  ]r^  (hhe]r_  (hh	e]r`  (hhe]ra  (jc  ]rb  (hh	e]rc  (hh	eeee]rd  (hheeejW  jW  jW  jW  jW  jW  jW  ]re  (jF  ]rf  (jH  ]rg  (jJ  ]rh  (hh	e]ri  (hhe]rj  (hjN  e]rk  (j^  ]rl  (hhe]rm  (hh	e]rn  (hhe]ro  (jc  ]rp  (hh	e]rq  (hh	eeee]rr  (hheeeje  je  je  je  je  ]rs  (jF  ]rt  (jH  ]ru  (jJ  ]rv  (hh	e]rw  (hhe]rx  (hjN  e]ry  (j^  ]rz  (hhe]r{  (hh	e]r|  (hhe]r}  (jc  ]r~  (hh	e]r  (hh	eeee]r�  (hheeejs  js  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r   (jH  ]r  (jJ  ]r  (hh	e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r	  (jc  ]r
  (hh	e]r  (hh	eeee]r  (hheeej�  j�  j�  j�  j�  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh	e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheeej  j  j  j  j  j  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh	e]r  (hhe]r   (hjN  e]r!  (j^  ]r"  (hhe]r#  (hh	e]r$  (hhe]r%  (jc  ]r&  (hh	e]r'  (hh	eeee]r(  (hheeej  j  j  j  j  j  ]r)  (jF  ]r*  (jH  ]r+  (jJ  ]r,  (hh	e]r-  (hhe]r.  (hjN  e]r/  (j^  ]r0  (hhe]r1  (hh	e]r2  (hhe]r3  (jc  ]r4  (hh	e]r5  (hh	eeee]r6  (hheeej)  ]r7  (jF  ]r8  (jH  ]r9  (jJ  ]r:  (hh	e]r;  (hhe]r<  (hjN  e]r=  (j^  ]r>  (hhe]r?  (hh	e]r@  (hhe]rA  (jc  ]rB  (hh	e]rC  (hh	eeee]rD  (hheeej7  ]rE  (jF  ]rF  (jH  ]rG  (jJ  ]rH  (hh	e]rI  (hhe]rJ  (hjN  e]rK  (j^  ]rL  (hhe]rM  (hh	e]rN  (hhe]rO  (jc  ]rP  (hh	e]rQ  (hh	eeee]rR  (hheeejE  jE  jE  ]rS  (jF  ]rT  (jH  ]rU  (jJ  ]rV  (hh	e]rW  (hhe]rX  (hjN  e]rY  (j^  ]rZ  (hhe]r[  (hh	e]r\  (hhe]r]  (jc  ]r^  (hh	e]r_  (hh	eeee]r`  (hheeejS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  jS  ]ra  (jF  ]rb  (jH  ]rc  (jJ  ]rd  (hh	e]re  (hhe]rf  (hjN  e]rg  (j^  ]rh  (hhe]ri  (hh	e]rj  (hhe]rk  (jc  ]rl  (hh	e]rm  (hh	eeee]rn  (hheeeja  ja  ja  ja  ja  ]ro  (jF  ]rp  (jH  ]rq  (jJ  ]rr  (hh	e]rs  (hhe]rt  (hjN  e]ru  (j^  ]rv  (hhe]rw  (hh	e]rx  (hhe]ry  (jc  ]rz  (hh	e]r{  (hh	eeee]r|  (hheeejo  jo  ]r}  (jF  ]r~  (jH  ]r  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej}  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r   (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheeej�  ]r	  (jF  ]r
  (jH  ]r  (jJ  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheeej	  j	  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r   (hhe]r!  (jc  ]r"  (hh	e]r#  (hh	eeee]r$  (hheee]r%  (jF  ]r&  (jH  ]r'  (jJ  ]r(  (hh"e]r)  (hhe]r*  (hjN  e]r+  (j^  ]r,  (hhe]r-  (hh	e]r.  (hhe]r/  (jc  ]r0  (hh	e]r1  (hh	eeee]r2  (hheeej%  j%  ]r3  (jF  ]r4  (jH  ]r5  (jJ  ]r6  (hh	e]r7  (hhe]r8  (hjN  e]r9  (j^  ]r:  (hhe]r;  (hh	e]r<  (hhe]r=  (jc  ]r>  (hh	e]r?  (hh	eeee]r@  (hheee]rA  (jF  ]rB  (jH  ]rC  (jJ  ]rD  (hh	e]rE  (hhe]rF  (hjN  e]rG  (j^  ]rH  (hhe]rI  (hh	e]rJ  (hhe]rK  (jc  ]rL  (hh	e]rM  (hh	eeee]rN  (hheeejA  jA  jA  jA  ]rO  (jF  ]rP  (jH  ]rQ  (jJ  ]rR  (hh	e]rS  (hhe]rT  (hjN  e]rU  (j^  ]rV  (hhe]rW  (hh	e]rX  (hhe]rY  (jc  ]rZ  (hh	e]r[  (hh	eeee]r\  (hheeejO  ]r]  (jF  ]r^  (jH  ]r_  (jJ  ]r`  (hh	e]ra  (hhe]rb  (hjN  e]rc  (j^  ]rd  (hhe]re  (hh	e]rf  (hhe]rg  (jc  ]rh  (hh	e]ri  (hh	eeee]rj  (hheeej]  ]rk  (jF  ]rl  (jH  ]rm  (jJ  ]rn  (hh	e]ro  (hhe]rp  (hjN  e]rq  (j^  ]rr  (hhe]rs  (hh	e]rt  (hhe]ru  (jc  ]rv  (hh	e]rw  (hh	eeee]rx  (hheeejk  jk  jk  jk  jk  jk  ]ry  (jF  ]rz  (jH  ]r{  (jJ  ]r|  (hh	e]r}  (hhe]r~  (hjN  e]r  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeejy  jy  jy  jy  jy  jy  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r   (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheeej�  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r	  (hhe]r
  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheeej  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r   (hheee]r!  (jF  ]r"  (jH  ]r#  (jJ  ]r$  (hh"e]r%  (hhe]r&  (hjN  e]r'  (j^  ]r(  (hhe]r)  (hh	e]r*  (hhe]r+  (jc  ]r,  (hh	e]r-  (hh	eeee]r.  (hheeej!  j!  j!  ]r/  (jF  ]r0  (jH  ]r1  (jJ  ]r2  (hh	e]r3  (hhe]r4  (hjN  e]r5  (j^  ]r6  (hhe]r7  (hh	e]r8  (hhe]r9  (jc  ]r:  (hh	e]r;  (hh	eeee]r<  (hheeej/  j/  ]r=  (jF  ]r>  (jH  ]r?  (jJ  ]r@  (hh	e]rA  (hhe]rB  (hjN  e]rC  (j^  ]rD  (hhe]rE  (hh	e]rF  (hhe]rG  (jc  ]rH  (hh	e]rI  (hh	eeee]rJ  (hheee]rK  (jF  ]rL  (jH  ]rM  (jJ  ]rN  (hh	e]rO  (hhe]rP  (hjN  e]rQ  (j^  ]rR  (hhe]rS  (hh	e]rT  (hhe]rU  (jc  ]rV  (hh	e]rW  (hh	eeee]rX  (hheeejK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  ]rY  (jF  ]rZ  (jH  ]r[  (jJ  ]r\  (hh	e]r]  (hhe]r^  (hjN  e]r_  (j^  ]r`  (hhe]ra  (hh	e]rb  (hhe]rc  (jc  ]rd  (hh	e]re  (hh	eeee]rf  (hheee]rg  (jF  ]rh  (jH  ]ri  (jJ  ]rj  (hh	e]rk  (hhe]rl  (hjN  e]rm  (j^  ]rn  (hhe]ro  (hh	e]rp  (hhe]rq  (jc  ]rr  (hh	e]rs  (hh	eeee]rt  (hheee]ru  (jF  ]rv  (jH  ]rw  (jJ  ]rx  (hh	e]ry  (hhe]rz  (hjN  e]r{  (j^  ]r|  (hhe]r}  (hh	e]r~  (hhe]r  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeeju  ju  ju  ju  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh	e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  ]r�  (jF  ]r�  (jH  ]r�  (jJ  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j^  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (jc  ]r�  (hh	e]r�  (hh	eeee]r   (hheeej�  j�  j�  j�  j�  j�  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r	  (hh	e]r
  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheeej  ]r  (jF  ]r  (jH  ]r  (jJ  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (j^  ]r  (hhe]r  (hh	e]r  (hhe]r  (jc  ]r  (hh	e]r  (hh	eeee]r  (hheeej  j  j  j  j  j  j  j  ]r  (jF  ]r  (jH  ]r  (jJ  ]r   (hh"e]r!  (hhe]r"  (hjN  e]r#  (j^  ]r$  (hhe]r%  (hh	e]r&  (hhe]r'  (jc  ]r(  (hh	e]r)  (hh	eeee]r*  (hheeej  j  j  j  j  j  j  ]r+  (jF  ]r,  (jH  ]r-  (jJ  ]r.  (hh"e]r/  (hhe]r0  (hjN  e]r1  (j^  ]r2  (hhe]r3  (hh	e]r4  (hhe]r5  (jc  ]r6  (hh	e]r7  (hh	eeee]r8  (hheeej+  j+  j+  j+  j+  j+  j+  ]r9  (jF  ]r:  (jH  ]r;  (jJ  ]r<  (hh"e]r=  (hhe]r>  (hjN  e]r?  (j^  ]r@  (hhe]rA  (hh	e]rB  (hhe]rC  (jc  ]rD  (hh	e]rE  (hh	eeee]rF  (hheeej9  j9  j9  j9  j9  j9  ]rG  (jF  ]rH  (jH  ]rI  (jJ  ]rJ  (hh"e]rK  (hhe]rL  (hjN  e]rM  (j^  ]rN  (hhe]rO  (hh	e]rP  (hhe]rQ  (jc  ]rR  (hh	e]rS  (hh	eeee]rT  (hheee]rU  (jF  ]rV  (jH  ]rW  (jJ  ]rX  (hh"e]rY  (hhe]rZ  (hjN  e]r[  (j^  ]r\  (hhe]r]  (hh	e]r^  (hhe]r_  (jc  ]r`  (hh	e]ra  (hh	eeee]rb  (hheeejU  jU  jU  jU  jU  jU  jU  jU  ]rc  (jF  ]rd  (jH  ]re  (jJ  ]rf  (hh"e]rg  (hhe]rh  (hjN  e]ri  (j^  ]rj  (hhe]rk  (hh	e]rl  (hhe]rm  (jc  ]rn  (hh	e]ro  (hh	eeee]rp  (hheeejc  jc  jc  e(]rq  (X   Normrr  ]rs  (X   Oblrt  ]ru  (X   Movedrv  ]rw  (hh"e]rx  (hhe]ry  (hjN  e]rz  (X   Movedr{  ]r|  (hhe]r}  (hh	e]r~  (hhe]r  (X	   Next-Mover�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeejq  ]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  ]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  ]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  ]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r   (hh	eeee]r  (hheeej�  j�  j�  j�  j�  j�  ]r  (jr  ]r  (jt  ]r  (jv  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (j{  ]r	  (hhe]r
  (hh	e]r  (hhe]r  (j�  ]r  (hh	e]r  (hh	eeee]r  (hheeej  j  j  j  j  ]r  (jr  ]r  (jt  ]r  (jv  ]r  (hh"e]r  (hhe]r  (hjN  e]r  (j{  ]r  (hhe]r  (hh	e]r  (hhe]r  (j�  ]r  (hh	e]r  (hh	eeee]r  (hheee]r  (jr  ]r  (jt  ]r   (jv  ]r!  (hh"e]r"  (hhe]r#  (hjN  e]r$  (j{  ]r%  (hhe]r&  (hh	e]r'  (hhe]r(  (j�  ]r)  (hh	e]r*  (hh	eeee]r+  (hheee]r,  (jr  ]r-  (jt  ]r.  (jv  ]r/  (hh"e]r0  (hhe]r1  (hjN  e]r2  (j{  ]r3  (hhe]r4  (hh	e]r5  (hhe]r6  (j�  ]r7  (hh	e]r8  (hh	eeee]r9  (hheee]r:  (jr  ]r;  (jt  ]r<  (jv  ]r=  (hh"e]r>  (hhe]r?  (hjN  e]r@  (j{  ]rA  (hhe]rB  (hh	e]rC  (hhe]rD  (j�  ]rE  (hh	e]rF  (hh	eeee]rG  (hheeej:  j:  j:  ]rH  (jr  ]rI  (jt  ]rJ  (jv  ]rK  (hh"e]rL  (hhe]rM  (hjN  e]rN  (j{  ]rO  (hhe]rP  (hh	e]rQ  (hhe]rR  (j�  ]rS  (hh	e]rT  (hh	eeee]rU  (hheee]rV  (jr  ]rW  (jt  ]rX  (jv  ]rY  (hh"e]rZ  (hhe]r[  (hjN  e]r\  (j{  ]r]  (hhe]r^  (hh	e]r_  (hhe]r`  (j�  ]ra  (hh	e]rb  (hh	eeee]rc  (hheee]rd  (jr  ]re  (jt  ]rf  (jv  ]rg  (hh"e]rh  (hhe]ri  (hjN  e]rj  (j{  ]rk  (hhe]rl  (hh	e]rm  (hhe]rn  (j�  ]ro  (hh	e]rp  (hh	eeee]rq  (hheeejd  jd  jd  ]rr  (jr  ]rs  (jt  ]rt  (jv  ]ru  (hh"e]rv  (hhe]rw  (hjN  e]rx  (j{  ]ry  (hhe]rz  (hh	e]r{  (hhe]r|  (j�  ]r}  (hh	e]r~  (hh	eeee]r  (hheeejr  jr  jr  jr  jr  jr  jr  jr  jr  jr  jr  jr  jr  ]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  ]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  ]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  ]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheee]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  ]r�  (jr  ]r�  (jt  ]r�  (jv  ]r�  (hh"e]r�  (hhe]r�  (hjN  e]r�  (j{  ]r�  (hhe]r�  (hh	e]r�  (hhe]r�  (j�  ]r�  (hh	e]r�  (hh	eeee]r�  (hheeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (jr  ]r�  (jt  ]r    (jv  ]r   (hh"e]r   (hhe]r   (hjN  e]r   (j{  ]r   (hhe]r   (hh	e]r   (hhe]r   (j�  ]r	   (hh	e]r
   (hh	eeee]r   (hheee]r   (jr  ]r   (jt  ]r   (jv  ]r   (hh"e]r   (hh	e]r   (hjN  e]r   (j{  ]r   (hhe]r   (hh	e]r   (hhe]r   (j�  ]r   (hh	e]r   (hh	eeee]r   (hheeej   ]r   (jr  ]r   (jt  ]r   (jv  ]r   (hh"e]r   (hh	e]r   (hjN  e]r    (j{  ]r!   (hhe]r"   (hh	e]r#   (hhe]r$   (j�  ]r%   (hh	e]r&   (hh	eeee]r'   (hheeej   j   j   j   ]r(   (jr  ]r)   (jt  ]r*   (jv  ]r+   (hh"e]r,   (hh	e]r-   (hjN  e]r.   (j{  ]r/   (hhe]r0   (hh	e]r1   (hhe]r2   (j�  ]r3   (hh	e]r4   (hh	eeee]r5   (hheeej(   j(   ]r6   (jr  ]r7   (jt  ]r8   (jv  ]r9   (hh"e]r:   (hh	e]r;   (hjN  e]r<   (j{  ]r=   (hhe]r>   (hh	e]r?   (hhe]r@   (j�  ]rA   (hh	e]rB   (hh	eeee]rC   (hheee]rD   (jr  ]rE   (jt  ]rF   (jv  ]rG   (hh"e]rH   (hh	e]rI   (hjN  e]rJ   (j{  ]rK   (hhe]rL   (hh	e]rM   (hhe]rN   (j�  ]rO   (hh	e]rP   (hh	eeee]rQ   (hheee]rR   (jr  ]rS   (jt  ]rT   (jv  ]rU   (hh"e]rV   (hh	e]rW   (hjN  e]rX   (j{  ]rY   (hhe]rZ   (hh	e]r[   (hhe]r\   (j�  ]r]   (hh	e]r^   (hh	eeee]r_   (hheeejR   jR   jR   ]r`   (jr  ]ra   (jt  ]rb   (jv  ]rc   (hh"e]rd   (hh	e]re   (hjN  e]rf   (j{  ]rg   (hhe]rh   (hh	e]ri   (hhe]rj   (j�  ]rk   (hh	e]rl   (hh	eeee]rm   (hheee]rn   (jr  ]ro   (jt  ]rp   (jv  ]rq   (hh"e]rr   (hh	e]rs   (hjN  e]rt   (j{  ]ru   (hhe]rv   (hh	e]rw   (hhe]rx   (j�  ]ry   (hh	e]rz   (hh	eeee]r{   (hheee]r|   (jr  ]r}   (jt  ]r~   (jv  ]r   (hh"e]r�   (hh	e]r�   (hjN  e]r�   (j{  ]r�   (hhe]r�   (hh	e]r�   (hhe]r�   (j�  ]r�   (hh	e]r�   (hh	eeee]r�   (hheeej|   j|   ]r�   (jr  ]r�   (jt  ]r�   (jv  ]r�   (hh"e]r�   (hh	e]r�   (hjN  e]r�   (j{  ]r�   (hhe]r�   (hh	e]r�   (hhe]r�   (j�  ]r�   (hh	e]r�   (hh	eeee]r�   (hheeej�   j�   j�   j�   j�   j�   j�   j�   j�   j�   j�   j�   j�   j�   j�   ]r�   (jr  ]r�   (jt  ]r�   (jv  ]r�   (hh"e]r�   (hh	e]r�   (hjN  e]r�   (j{  ]r�   (hhe]r�   (hh	e]r�   (hhe]r�   (j�  ]r�   (hh	e]r�   (hh	eeee]r�   (hheeej�   j�   j�   ]r�   (jr  ]r�   (jt  ]r�   (jv  ]r�   (hh"e]r�   (hh	e]r�   (hjN  e]r�   (j{  ]r�   (hhe]r�   (hh	e]r�   (hhe]r�   (j�  ]r�   (hh	e]r�   (hh	eeee]r�   (hheeej�   j�   j�   j�   j�   ]r�   (jr  ]r�   (jt  ]r�   (jv  ]r�   (hh"e]r�   (hh	e]r�   (hjN  e]r�   (j{  ]r�   (hhe]r�   (hh	e]r�   (hhe]r�   (j�  ]r�   (hh	e]r�   (hh	eeee]r�   (hheeej�   j�   j�   j�   j�   ]r�   (jr  ]r�   (jt  ]r�   (jv  ]r�   (hh"e]r�   (hh	e]r�   (hjN  e]r�   (j{  ]r�   (hhe]r�   (hh	e]r�   (hhe]r�   (j�  ]r�   (hh	e]r�   (hh	eeee]r�   (hheeej�   j�   j�   j�   j�   j�   ]r�   (jr  ]r�   (jt  ]r�   (jv  ]r�   (hh"e]r�   (hh	e]r�   (hjN  e]r�   (j{  ]r�   (hhe]r�   (hh	e]r�   (hhe]r�   (j�  ]r�   (hh	e]r�   (hh	eeee]r�   (hheeej�   j�   ]r�   (jr  ]r�   (jt  ]r�   (jv  ]r�   (hh"e]r�   (hh	e]r�   (hjN  e]r�   (j{  ]r�   (hhe]r�   (hh	e]r�   (hhe]r�   (j�  ]r�   (hh	e]r�   (hh	eeee]r�   (hheee]r�   (jr  ]r�   (jt  ]r�   (jv  ]r�   (hh"e]r�   (hh	e]r�   (hjN  e]r�   (j{  ]r�   (hhe]r�   (hh	e]r�   (hhe]r�   (j�  ]r�   (hh	e]r�   (hh	eeee]r�   (hheeej�   j�   j�   ]r�   (jr  ]r�   (jt  ]r�   (jv  ]r�   (hh"e]r�   (hh	e]r�   (hjN  e]r !  (j{  ]r!  (hhe]r!  (hh	e]r!  (hhe]r!  (j�  ]r!  (hh	e]r!  (hh	eeee]r!  (hheeej�   j�   j�   ]r!  (jr  ]r	!  (jt  ]r
!  (jv  ]r!  (hh"e]r!  (hh	e]r!  (hjN  e]r!  (j{  ]r!  (hhe]r!  (hh	e]r!  (hhe]r!  (j�  ]r!  (hh	e]r!  (hh	eeee]r!  (hheeej!  j!  ]r!  (jr  ]r!  (jt  ]r!  (jv  ]r!  (hh"e]r!  (hh	e]r!  (hjN  e]r!  (j{  ]r!  (hhe]r!  (hh	e]r!  (hhe]r !  (j�  ]r!!  (hh	e]r"!  (hh	eeee]r#!  (hheeej!  j!  ]r$!  (jr  ]r%!  (jt  ]r&!  (jv  ]r'!  (hh"e]r(!  (hh	e]r)!  (hjN  e]r*!  (j{  ]r+!  (hhe]r,!  (hh	e]r-!  (hhe]r.!  (j�  ]r/!  (hh	e]r0!  (hh	eeee]r1!  (hheeej$!  j$!  ]r2!  (jr  ]r3!  (jt  ]r4!  (jv  ]r5!  (hh"e]r6!  (hh	e]r7!  (hjN  e]r8!  (j{  ]r9!  (hhe]r:!  (hh	e]r;!  (hhe]r<!  (j�  ]r=!  (hh	e]r>!  (hh	eeee]r?!  (hheeej2!  j2!  j2!  j2!  j2!  j2!  j2!  ]r@!  (jr  ]rA!  (jt  ]rB!  (jv  ]rC!  (hh"e]rD!  (hh	e]rE!  (hjN  e]rF!  (j{  ]rG!  (hhe]rH!  (hh	e]rI!  (hhe]rJ!  (j�  ]rK!  (hh	e]rL!  (hh	eeee]rM!  (hheee]rN!  (jr  ]rO!  (jt  ]rP!  (jv  ]rQ!  (hh"e]rR!  (hh	e]rS!  (hjN  e]rT!  (j{  ]rU!  (hhe]rV!  (hh	e]rW!  (hhe]rX!  (j�  ]rY!  (hh	e]rZ!  (hh	eeee]r[!  (hheeejN!  jN!  jN!  ]r\!  (jr  ]r]!  (jt  ]r^!  (jv  ]r_!  (hh"e]r`!  (hh	e]ra!  (hjN  e]rb!  (j{  ]rc!  (hhe]rd!  (hh	e]re!  (hhe]rf!  (j�  ]rg!  (hh	e]rh!  (hh	eeee]ri!  (hheeej\!  ]rj!  (jr  ]rk!  (jt  ]rl!  (jv  ]rm!  (hh"e]rn!  (hh	e]ro!  (hjN  e]rp!  (j{  ]rq!  (hhe]rr!  (hh	e]rs!  (hhe]rt!  (j�  ]ru!  (hh	e]rv!  (hh	eeee]rw!  (hheeejj!  jj!  jj!  jj!  jj!  ]rx!  (jr  ]ry!  (jt  ]rz!  (jv  ]r{!  (hh"e]r|!  (hh	e]r}!  (hjN  e]r~!  (j{  ]r!  (hhe]r�!  (hh	e]r�!  (hhe]r�!  (j�  ]r�!  (hh	e]r�!  (hh	eeee]r�!  (hheee]r�!  (jr  ]r�!  (jt  ]r�!  (jv  ]r�!  (hh"e]r�!  (hh	e]r�!  (hjN  e]r�!  (j{  ]r�!  (hhe]r�!  (hh	e]r�!  (hhe]r�!  (j�  ]r�!  (hh	e]r�!  (hh	eeee]r�!  (hheeej�!  j�!  j�!  j�!  j�!  j�!  j�!  j�!  ]r�!  (jr  ]r�!  (jt  ]r�!  (jv  ]r�!  (hh"e]r�!  (hhe]r�!  (hjN  e]r�!  (j{  ]r�!  (hhe]r�!  (hh	e]r�!  (hhe]r�!  (j�  ]r�!  (hh	e]r�!  (hh	eeee]r�!  (hheeej�!  j�!  j�!  j�!  j�!  ]r�!  (jr  ]r�!  (jt  ]r�!  (jv  ]r�!  (hh"e]r�!  (hhe]r�!  (hjN  e]r�!  (j{  ]r�!  (hhe]r�!  (hh	e]r�!  (hhe]r�!  (j�  ]r�!  (hh	e]r�!  (hh	eeee]r�!  (hheeej�!  j�!  j�!  j�!  ]r�!  (jr  ]r�!  (jt  ]r�!  (jv  ]r�!  (hh"e]r�!  (hhe]r�!  (hjN  e]r�!  (j{  ]r�!  (hhe]r�!  (hh	e]r�!  (hhe]r�!  (j�  ]r�!  (hh	e]r�!  (hh	eeee]r�!  (hheee]r�!  (jr  ]r�!  (jt  ]r�!  (jv  ]r�!  (hh"e]r�!  (hhe]r�!  (hjN  e]r�!  (j{  ]r�!  (hhe]r�!  (hh	e]r�!  (hhe]r�!  (j�  ]r�!  (hh	e]r�!  (hh	eeee]r�!  (hheee]r�!  (jr  ]r�!  (jt  ]r�!  (jv  ]r�!  (hh"e]r�!  (hhe]r�!  (hjN  e]r�!  (j{  ]r�!  (hhe]r�!  (hh	e]r�!  (hhe]r�!  (j�  ]r�!  (hh	e]r�!  (hh	eeee]r�!  (hheeej�!  ]r�!  (jr  ]r�!  (jt  ]r�!  (jv  ]r�!  (hh"e]r�!  (hhe]r�!  (hjN  e]r�!  (j{  ]r�!  (hhe]r�!  (hh	e]r�!  (hhe]r�!  (j�  ]r�!  (hh	e]r�!  (hh	eeee]r�!  (hheeej�!  j�!  j�!  j�!  j�!  ]r�!  (jr  ]r�!  (jt  ]r�!  (jv  ]r�!  (hh"e]r�!  (hhe]r�!  (hjN  e]r�!  (j{  ]r�!  (hhe]r�!  (hh	e]r�!  (hhe]r�!  (j�  ]r�!  (hh	e]r�!  (hh	eeee]r�!  (hheee]r�!  (jr  ]r�!  (jt  ]r�!  (jv  ]r�!  (hh"e]r�!  (hh	e]r�!  (hjN  e]r�!  (j{  ]r�!  (hhe]r�!  (hh	e]r�!  (hhe]r "  (j�  ]r"  (hh	e]r"  (hh	eeee]r"  (hheee]r"  (jr  ]r"  (jt  ]r"  (jv  ]r"  (hh"e]r"  (hh	e]r	"  (hjN  e]r
"  (j{  ]r"  (hhe]r"  (hh	e]r"  (hhe]r"  (j�  ]r"  (hh	e]r"  (hh	eeee]r"  (hheeej"  j"  j"  ]r"  (jr  ]r"  (jt  ]r"  (jv  ]r"  (hh"e]r"  (hh	e]r"  (hjN  e]r"  (j{  ]r"  (hhe]r"  (hh	e]r"  (hhe]r"  (j�  ]r"  (hh	e]r"  (hh	eeee]r"  (hheeej"  ]r "  (jr  ]r!"  (jt  ]r""  (jv  ]r#"  (hh"e]r$"  (hh	e]r%"  (hjN  e]r&"  (j{  ]r'"  (hhe]r("  (hh	e]r)"  (hhe]r*"  (j�  ]r+"  (hh	e]r,"  (hh	eeee]r-"  (hheeej "  ]r."  (jr  ]r/"  (jt  ]r0"  (jv  ]r1"  (hh"e]r2"  (hh	e]r3"  (hjN  e]r4"  (j{  ]r5"  (hhe]r6"  (hh	e]r7"  (hhe]r8"  (j�  ]r9"  (hh	e]r:"  (hh	eeee]r;"  (hheeej."  j."  j."  j."  ]r<"  (jr  ]r="  (jt  ]r>"  (jv  ]r?"  (hh"e]r@"  (hh	e]rA"  (hjN  e]rB"  (j{  ]rC"  (hhe]rD"  (hh	e]rE"  (hhe]rF"  (j�  ]rG"  (hh	e]rH"  (hh	eeee]rI"  (hheeej<"  j<"  ]rJ"  (jr  ]rK"  (jt  ]rL"  (jv  ]rM"  (hh"e]rN"  (hh	e]rO"  (hjN  e]rP"  (j{  ]rQ"  (hhe]rR"  (hh	e]rS"  (hhe]rT"  (j�  ]rU"  (hh	e]rV"  (hh	eeee]rW"  (hheeejJ"  jJ"  ]rX"  (jr  ]rY"  (jt  ]rZ"  (jv  ]r["  (hh"e]r\"  (hh	e]r]"  (hjN  e]r^"  (j{  ]r_"  (hhe]r`"  (hh	e]ra"  (hhe]rb"  (j�  ]rc"  (hh	e]rd"  (hh	eeee]re"  (hheeejX"  jX"  jX"  jX"  jX"  jX"  jX"  jX"  jX"  jX"  ]rf"  (jr  ]rg"  (jt  ]rh"  (jv  ]ri"  (hh"e]rj"  (hh	e]rk"  (hjN  e]rl"  (j{  ]rm"  (hhe]rn"  (hh	e]ro"  (hhe]rp"  (j�  ]rq"  (hh	e]rr"  (hh	eeee]rs"  (hheee]rt"  (jr  ]ru"  (jt  ]rv"  (jv  ]rw"  (hh"e]rx"  (hh	e]ry"  (hjN  e]rz"  (j{  ]r{"  (hhe]r|"  (hh	e]r}"  (hhe]r~"  (j�  ]r"  (hh	e]r�"  (hh	eeee]r�"  (hheeejt"  jt"  jt"  ]r�"  (jr  ]r�"  (jt  ]r�"  (jv  ]r�"  (hh"e]r�"  (hhe]r�"  (hjN  e]r�"  (j{  ]r�"  (hhe]r�"  (hh	e]r�"  (hhe]r�"  (j�  ]r�"  (hh	e]r�"  (hh	eeee]r�"  (hheeej�"  j�"  j�"  j�"  j�"  j�"  j�"  j�"  j�"  j�"  j�"  j�"  j�"  j�"  j�"  ]r�"  (jr  ]r�"  (jt  ]r�"  (jv  ]r�"  (hh"e]r�"  (hhe]r�"  (hjN  e]r�"  (j{  ]r�"  (hhe]r�"  (hh	e]r�"  (hhe]r�"  (j�  ]r�"  (hh	e]r�"  (hh	eeee]r�"  (hheeej�"  j�"  ]r�"  (jr  ]r�"  (jt  ]r�"  (jv  ]r�"  (hh"e]r�"  (hhe]r�"  (hjN  e]r�"  (j{  ]r�"  (hhe]r�"  (hh	e]r�"  (hhe]r�"  (j�  ]r�"  (hh	e]r�"  (hh	eeee]r�"  (hheeej�"  j�"  j�"  j�"  j�"  j�"  j�"  j�"  j�"  ]r�"  (jr  ]r�"  (jt  ]r�"  (jv  ]r�"  (hh"e]r�"  (hhe]r�"  (hjN  e]r�"  (j{  ]r�"  (hhe]r�"  (hh	e]r�"  (hhe]r�"  (j�  ]r�"  (hh	e]r�"  (hh	eeee]r�"  (hheee]r�"  (jr  ]r�"  (jt  ]r�"  (jv  ]r�"  (hh"e]r�"  (hhe]r�"  (hjN  e]r�"  (j{  ]r�"  (hhe]r�"  (hh	e]r�"  (hhe]r�"  (j�  ]r�"  (hh	e]r�"  (hh	eeee]r�"  (hheeej�"  j�"  j�"  ]r�"  (jr  ]r�"  (jt  ]r�"  (jv  ]r�"  (hh"e]r�"  (hhe]r�"  (hjN  e]r�"  (j{  ]r�"  (hhe]r�"  (hh	e]r�"  (hhe]r�"  (j�  ]r�"  (hh	e]r�"  (hh	eeee]r�"  (hheeej�"  j�"  j�"  j�"  j�"  j�"  ]r�"  (jr  ]r�"  (jt  ]r�"  (jv  ]r�"  (hh"e]r�"  (hhe]r�"  (hjN  e]r�"  (j{  ]r�"  (hhe]r�"  (hh	e]r�"  (hhe]r�"  (j�  ]r�"  (hh	e]r�"  (hh	eeee]r�"  (hheeej�"  ]r�"  (jr  ]r�"  (jt  ]r�"  (jv  ]r�"  (hh"e]r�"  (hh	e]r�"  (hjN  e]r�"  (j{  ]r�"  (hhe]r�"  (hh	e]r�"  (hhe]r�"  (j�  ]r�"  (hh	e]r�"  (hh	eeee]r�"  (hheeej�"  j�"  ]r�"  (jr  ]r�"  (jt  ]r�"  (jv  ]r�"  (hh"e]r�"  (hh	e]r�"  (hjN  e]r�"  (j{  ]r�"  (hhe]r�"  (hh	e]r�"  (hhe]r�"  (j�  ]r�"  (hh	e]r�"  (hh	eeee]r�"  (hheeej�"  j�"  j�"  j�"  ]r #  (jr  ]r#  (jt  ]r#  (jv  ]r#  (hh"e]r#  (hh	e]r#  (hjN  e]r#  (j{  ]r#  (hhe]r#  (hh	e]r	#  (hhe]r
#  (j�  ]r#  (hh	e]r#  (hh	eeee]r#  (hheeej #  ]r#  (jr  ]r#  (jt  ]r#  (jv  ]r#  (hh"e]r#  (hh	e]r#  (hjN  e]r#  (j{  ]r#  (hhe]r#  (hh	e]r#  (hhe]r#  (j�  ]r#  (hh	e]r#  (hh	eeee]r#  (hheeej#  j#  j#  j#  j#  j#  j#  j#  j#  j#  j#  j#  ]r#  (jr  ]r#  (jt  ]r#  (jv  ]r#  (hh"e]r #  (hh	e]r!#  (hjN  e]r"#  (j{  ]r##  (hhe]r$#  (hh	e]r%#  (hhe]r&#  (j�  ]r'#  (hh	e]r(#  (hh	eeee]r)#  (hheee]r*#  (jr  ]r+#  (jt  ]r,#  (jv  ]r-#  (hh"e]r.#  (hh	e]r/#  (hjN  e]r0#  (j{  ]r1#  (hhe]r2#  (hh	e]r3#  (hhe]r4#  (j�  ]r5#  (hh	e]r6#  (hh	eeee]r7#  (hheeej*#  j*#  j*#  j*#  j*#  j*#  j*#  ]r8#  (jr  ]r9#  (jt  ]r:#  (jv  ]r;#  (hh"e]r<#  (hh	e]r=#  (hjN  e]r>#  (j{  ]r?#  (hhe]r@#  (hh	e]rA#  (hhe]rB#  (j�  ]rC#  (hh	e]rD#  (hh	eeee]rE#  (hheee]rF#  (jr  ]rG#  (jt  ]rH#  (jv  ]rI#  (hh"e]rJ#  (hh	e]rK#  (hjN  e]rL#  (j{  ]rM#  (hhe]rN#  (hh	e]rO#  (hhe]rP#  (j�  ]rQ#  (hh	e]rR#  (hh	eeee]rS#  (hheeejF#  jF#  jF#  jF#  jF#  jF#  jF#  jF#  jF#  jF#  ]rT#  (jr  ]rU#  (jt  ]rV#  (jv  ]rW#  (hh"e]rX#  (hh	e]rY#  (hjN  e]rZ#  (j{  ]r[#  (hhe]r\#  (hh	e]r]#  (hhe]r^#  (j�  ]r_#  (hh	e]r`#  (hh	eeee]ra#  (hheeejT#  ]rb#  (jr  ]rc#  (jt  ]rd#  (jv  ]re#  (hh"e]rf#  (hh	e]rg#  (hjN  e]rh#  (j{  ]ri#  (hhe]rj#  (hh	e]rk#  (hhe]rl#  (j�  ]rm#  (hh	e]rn#  (hh	eeee]ro#  (hheeejb#  jb#  jb#  jb#  jb#  jb#  ]rp#  (jr  ]rq#  (jt  ]rr#  (jv  ]rs#  (hh"e]rt#  (hh	e]ru#  (hjN  e]rv#  (j{  ]rw#  (hhe]rx#  (hh	e]ry#  (hhe]rz#  (j�  ]r{#  (hh	e]r|#  (hh	eeee]r}#  (hheeejp#  jp#  jp#  jp#  jp#  jp#  jp#  jp#  jp#  jp#  jp#  jp#  jp#  jp#  jp#  jp#  ]r~#  (jr  ]r#  (jt  ]r�#  (jv  ]r�#  (hh"e]r�#  (hh	e]r�#  (hjN  e]r�#  (j{  ]r�#  (hhe]r�#  (hh	e]r�#  (hhe]r�#  (j�  ]r�#  (hh	e]r�#  (hh	eeee]r�#  (hheee]r�#  (jr  ]r�#  (jt  ]r�#  (jv  ]r�#  (hh"e]r�#  (hh	e]r�#  (hjN  e]r�#  (j{  ]r�#  (hhe]r�#  (hh	e]r�#  (hhe]r�#  (j�  ]r�#  (hh	e]r�#  (hh	eeee]r�#  (hheee]r�#  (jr  ]r�#  (jt  ]r�#  (jv  ]r�#  (hh"e]r�#  (hh	e]r�#  (hjN  e]r�#  (j{  ]r�#  (hhe]r�#  (hh	e]r�#  (hhe]r�#  (j�  ]r�#  (hh	e]r�#  (hh	eeee]r�#  (hheeej�#  j�#  ]r�#  (jr  ]r�#  (jt  ]r�#  (jv  ]r�#  (hh"e]r�#  (hhe]r�#  (hjN  e]r�#  (j{  ]r�#  (hhe]r�#  (hh	e]r�#  (hhe]r�#  (j�  ]r�#  (hh	e]r�#  (hh	eeee]r�#  (hheeej�#  j�#  j�#  ]r�#  (jr  ]r�#  (jt  ]r�#  (jv  ]r�#  (hh"e]r�#  (hhe]r�#  (hjN  e]r�#  (j{  ]r�#  (hhe]r�#  (hh	e]r�#  (hhe]r�#  (j�  ]r�#  (hh	e]r�#  (hh	eeee]r�#  (hheeej�#  j�#  ]r�#  (jr  ]r�#  (jt  ]r�#  (jv  ]r�#  (hh"e]r�#  (hhe]r�#  (hjN  e]r�#  (j{  ]r�#  (hhe]r�#  (hh	e]r�#  (hhe]r�#  (j�  ]r�#  (hh	e]r�#  (hh	eeee]r�#  (hheeej�#  j�#  j�#  j�#  j�#  j�#  j�#  ]r�#  (jr  ]r�#  (jt  ]r�#  (jv  ]r�#  (hh"e]r�#  (hhe]r�#  (hjN  e]r�#  (j{  ]r�#  (hhe]r�#  (hh	e]r�#  (hhe]r�#  (j�  ]r�#  (hh	e]r�#  (hh	eeee]r�#  (hheeej�#  j�#  j�#  j�#  j�#  j�#  j�#  j�#  j�#  j�#  ]r�#  (jr  ]r�#  (jt  ]r�#  (jv  ]r�#  (hh"e]r�#  (hhe]r�#  (hjN  e]r�#  (j{  ]r�#  (hhe]r�#  (hh	e]r�#  (hhe]r�#  (j�  ]r�#  (hh	e]r�#  (hh	eeee]r�#  (hheeej�#  j�#  j�#  j�#  j�#  ]r�#  (jr  ]r�#  (jt  ]r�#  (jv  ]r�#  (hh"e]r�#  (hhe]r�#  (hjN  e]r�#  (j{  ]r�#  (hhe]r�#  (hh	e]r�#  (hhe]r�#  (j�  ]r�#  (hh	e]r�#  (hh	eeee]r�#  (hheeej�#  j�#  j�#  j�#  j�#  j�#  j�#  j�#  j�#  j�#  j�#  j�#  ]r�#  (jr  ]r�#  (jt  ]r�#  (jv  ]r�#  (hh"e]r $  (hhe]r$  (hjN  e]r$  (j{  ]r$  (hhe]r$  (hh	e]r$  (hhe]r$  (j�  ]r$  (hh	e]r$  (hh	eeee]r	$  (hheeej�#  j�#  j�#  j�#  j�#  j�#  j�#  j�#  ]r
$  (jr  ]r$  (jt  ]r$  (jv  ]r$  (hh"e]r$  (hhe]r$  (hjN  e]r$  (j{  ]r$  (hhe]r$  (hh	e]r$  (hhe]r$  (j�  ]r$  (hh	e]r$  (hh	eeee]r$  (hheeej
$  j
$  ]r$  (jr  ]r$  (jt  ]r$  (jv  ]r$  (hh"e]r$  (hhe]r$  (hjN  e]r$  (j{  ]r$  (hhe]r $  (hh	e]r!$  (hhe]r"$  (j�  ]r#$  (hh	e]r$$  (hh	eeee]r%$  (hheeej$  j$  j$  ]r&$  (jr  ]r'$  (jt  ]r($  (jv  ]r)$  (hh"e]r*$  (hhe]r+$  (hjN  e]r,$  (j{  ]r-$  (hhe]r.$  (hh	e]r/$  (hhe]r0$  (j�  ]r1$  (hh	e]r2$  (hh	eeee]r3$  (hheeej&$  ]r4$  (jr  ]r5$  (jt  ]r6$  (jv  ]r7$  (hh"e]r8$  (hhe]r9$  (hjN  e]r:$  (j{  ]r;$  (hhe]r<$  (hh	e]r=$  (hhe]r>$  (j�  ]r?$  (hh	e]r@$  (hh	eeee]rA$  (hheeej4$  ]rB$  (jr  ]rC$  (jt  ]rD$  (jv  ]rE$  (hh"e]rF$  (hhe]rG$  (hjN  e]rH$  (j{  ]rI$  (hhe]rJ$  (hh	e]rK$  (hhe]rL$  (j�  ]rM$  (hh	e]rN$  (hh	eeee]rO$  (hheeejB$  jB$  jB$  ]rP$  (jr  ]rQ$  (jt  ]rR$  (jv  ]rS$  (hh"e]rT$  (hh	e]rU$  (hjN  e]rV$  (j{  ]rW$  (hhe]rX$  (hh	e]rY$  (hhe]rZ$  (j�  ]r[$  (hh	e]r\$  (hh	eeee]r]$  (hheee]r^$  (jr  ]r_$  (jt  ]r`$  (jv  ]ra$  (hh"e]rb$  (hhe]rc$  (hjN  e]rd$  (j{  ]re$  (hhe]rf$  (hh	e]rg$  (hhe]rh$  (j�  ]ri$  (hh	e]rj$  (hh	eeee]rk$  (hheeej^$  j^$  j^$  j^$  j^$  j^$  ]rl$  (jr  ]rm$  (jt  ]rn$  (jv  ]ro$  (hh"e]rp$  (hhe]rq$  (hjN  e]rr$  (j{  ]rs$  (hhe]rt$  (hh	e]ru$  (hhe]rv$  (j�  ]rw$  (hh	e]rx$  (hh	eeee]ry$  (hheeejl$  jl$  jl$  jl$  ]rz$  (jr  ]r{$  (jt  ]r|$  (jv  ]r}$  (hh"e]r~$  (hhe]r$  (hjN  e]r�$  (j{  ]r�$  (hhe]r�$  (hh	e]r�$  (hhe]r�$  (j�  ]r�$  (hh	e]r�$  (hh	eeee]r�$  (hheee]r�$  (jr  ]r�$  (jt  ]r�$  (jv  ]r�$  (hh"e]r�$  (hhe]r�$  (hjN  e]r�$  (j{  ]r�$  (hhe]r�$  (hh	e]r�$  (hhe]r�$  (j�  ]r�$  (hh	e]r�$  (hh	eeee]r�$  (hheeej�$  j�$  ]r�$  (jr  ]r�$  (jt  ]r�$  (jv  ]r�$  (hh"e]r�$  (hhe]r�$  (hjN  e]r�$  (j{  ]r�$  (hhe]r�$  (hh	e]r�$  (hhe]r�$  (j�  ]r�$  (hh	e]r�$  (hh	eeee]r�$  (hheeej�$  ]r�$  (jr  ]r�$  (jt  ]r�$  (jv  ]r�$  (hh"e]r�$  (hhe]r�$  (hjN  e]r�$  (j{  ]r�$  (hhe]r�$  (hh	e]r�$  (hhe]r�$  (j�  ]r�$  (hh	e]r�$  (hh	eeee]r�$  (hheeej�$  j�$  j�$  j�$  j�$  j�$  j�$  j�$  ]r�$  (jr  ]r�$  (jt  ]r�$  (jv  ]r�$  (hh"e]r�$  (hhe]r�$  (hjN  e]r�$  (j{  ]r�$  (hhe]r�$  (hh	e]r�$  (hhe]r�$  (j�  ]r�$  (hh	e]r�$  (hh	eeee]r�$  (hheeej�$  j�$  j�$  ]r�$  (jr  ]r�$  (jt  ]r�$  (jv  ]r�$  (hh"e]r�$  (hhe]r�$  (hjN  e]r�$  (j{  ]r�$  (hhe]r�$  (hh	e]r�$  (hhe]r�$  (j�  ]r�$  (hh	e]r�$  (hh	eeee]r�$  (hheeej�$  j�$  j�$  j�$  j�$  j�$  ]r�$  (jr  ]r�$  (jt  ]r�$  (jv  ]r�$  (hh"e]r�$  (hhe]r�$  (hjN  e]r�$  (j{  ]r�$  (hhe]r�$  (hh	e]r�$  (hhe]r�$  (j�  ]r�$  (hh	e]r�$  (hh	eeee]r�$  (hheeej�$  ]r�$  (jr  ]r�$  (jt  ]r�$  (jv  ]r�$  (hh"e]r�$  (hh	e]r�$  (hjN  e]r�$  (j{  ]r�$  (hhe]r�$  (hh	e]r�$  (hhe]r�$  (j�  ]r�$  (hh	e]r�$  (hh	eeee]r�$  (hheeej�$  j�$  j�$  ]r�$  (jr  ]r�$  (jt  ]r�$  (jv  ]r�$  (hh"e]r�$  (hh	e]r�$  (hjN  e]r�$  (j{  ]r�$  (hhe]r�$  (hh	e]r�$  (hhe]r�$  (j�  ]r�$  (hh	e]r�$  (hh	eeee]r�$  (hheee]r�$  (jr  ]r�$  (jt  ]r�$  (jv  ]r�$  (hh"e]r�$  (hh	e]r�$  (hjN  e]r�$  (j{  ]r�$  (hhe]r %  (hh	e]r%  (hhe]r%  (j�  ]r%  (hh	e]r%  (hh	eeee]r%  (hheeej�$  j�$  j�$  j�$  j�$  j�$  j�$  ]r%  (jr  ]r%  (jt  ]r%  (jv  ]r	%  (hh"e]r
%  (hh	e]r%  (hjN  e]r%  (j{  ]r%  (hhe]r%  (hh	e]r%  (hhe]r%  (j�  ]r%  (hh	e]r%  (hh	eeee]r%  (hheee]r%  (jr  ]r%  (jt  ]r%  (jv  ]r%  (hh"e]r%  (hh	e]r%  (hjN  e]r%  (j{  ]r%  (hhe]r%  (hh	e]r%  (hhe]r%  (j�  ]r%  (hh	e]r %  (hh	eeee]r!%  (hheee]r"%  (jr  ]r#%  (jt  ]r$%  (jv  ]r%%  (hh"e]r&%  (hh	e]r'%  (hjN  e]r(%  (j{  ]r)%  (hhe]r*%  (hh	e]r+%  (hhe]r,%  (j�  ]r-%  (hh	e]r.%  (hh	eeee]r/%  (hheee]r0%  (jr  ]r1%  (jt  ]r2%  (jv  ]r3%  (hh"e]r4%  (hh	e]r5%  (hjN  e]r6%  (j{  ]r7%  (hhe]r8%  (hh	e]r9%  (hhe]r:%  (j�  ]r;%  (hh	e]r<%  (hh	eeee]r=%  (hheeej0%  j0%  ]r>%  (jr  ]r?%  (jt  ]r@%  (jv  ]rA%  (hh"e]rB%  (hhe]rC%  (hjN  e]rD%  (j{  ]rE%  (hhe]rF%  (hh	e]rG%  (hhe]rH%  (j�  ]rI%  (hh	e]rJ%  (hh	eeee]rK%  (hheeej>%  ]rL%  (jr  ]rM%  (jt  ]rN%  (jv  ]rO%  (hh"e]rP%  (hhe]rQ%  (hjN  e]rR%  (j{  ]rS%  (hhe]rT%  (hh	e]rU%  (hhe]rV%  (j�  ]rW%  (hh	e]rX%  (hh	eeee]rY%  (hheeejL%  jL%  jL%  jL%  jL%  jL%  jL%  ]rZ%  (jr  ]r[%  (jt  ]r\%  (jv  ]r]%  (hh"e]r^%  (hhe]r_%  (hjN  e]r`%  (j{  ]ra%  (hhe]rb%  (hh	e]rc%  (hhe]rd%  (j�  ]re%  (hh	e]rf%  (hh	eeee]rg%  (hheee]rh%  (jr  ]ri%  (jt  ]rj%  (jv  ]rk%  (hh	e]rl%  (hhe]rm%  (hjN  e]rn%  (j{  ]ro%  (hhe]rp%  (hh	e]rq%  (hhe]rr%  (j�  ]rs%  (hh	e]rt%  (hh	eeee]ru%  (hheeejh%  jh%  ]rv%  (jr  ]rw%  (jt  ]rx%  (jv  ]ry%  (hh	e]rz%  (hhe]r{%  (hjN  e]r|%  (j{  ]r}%  (hhe]r~%  (hh	e]r%  (hhe]r�%  (j�  ]r�%  (hh	e]r�%  (hh	eeee]r�%  (hheeejv%  ]r�%  (jr  ]r�%  (jt  ]r�%  (jv  ]r�%  (hh	e]r�%  (hhe]r�%  (hjN  e]r�%  (j{  ]r�%  (hhe]r�%  (hh	e]r�%  (hhe]r�%  (j�  ]r�%  (hh	e]r�%  (hh	eeee]r�%  (hheeej�%  ]r�%  (jr  ]r�%  (jt  ]r�%  (jv  ]r�%  (hh	e]r�%  (hhe]r�%  (hjN  e]r�%  (j{  ]r�%  (hhe]r�%  (hh	e]r�%  (hhe]r�%  (j�  ]r�%  (hh	e]r�%  (hh	eeee]r�%  (hheeej�%  j�%  j�%  j�%  j�%  j�%  ]r�%  (jr  ]r�%  (jt  ]r�%  (jv  ]r�%  (hh	e]r�%  (hhe]r�%  (hjN  e]r�%  (j{  ]r�%  (hhe]r�%  (hh	e]r�%  (hhe]r�%  (j�  ]r�%  (hh	e]r�%  (hh	eeee]r�%  (hheeej�%  j�%  ]r�%  (jr  ]r�%  (jt  ]r�%  (jv  ]r�%  (hh	e]r�%  (hhe]r�%  (hjN  e]r�%  (j{  ]r�%  (hhe]r�%  (hh	e]r�%  (hhe]r�%  (j�  ]r�%  (hh	e]r�%  (hh	eeee]r�%  (hheeej�%  j�%  j�%  j�%  j�%  j�%  j�%  j�%  j�%  j�%  j�%  j�%  j�%  ]r�%  (jr  ]r�%  (jt  ]r�%  (jv  ]r�%  (hh"e]r�%  (hhe]r�%  (hjN  e]r�%  (j{  ]r�%  (hhe]r�%  (hh	e]r�%  (hhe]r�%  (j�  ]r�%  (hh	e]r�%  (hh	eeee]r�%  (hheeej�%  j�%  j�%  j�%  j�%  ]r�%  (jr  ]r�%  (jt  ]r�%  (jv  ]r�%  (hh"e]r�%  (hh	e]r�%  (hjN  e]r�%  (j{  ]r�%  (hhe]r�%  (hh	e]r�%  (hhe]r�%  (j�  ]r�%  (hh	e]r�%  (hh	eeee]r�%  (hheee]r�%  (jr  ]r�%  (jt  ]r�%  (jv  ]r�%  (hh"e]r�%  (hh	e]r�%  (hjN  e]r�%  (j{  ]r�%  (hhe]r�%  (hh	e]r�%  (hhe]r�%  (j�  ]r�%  (hh	e]r�%  (hh	eeee]r�%  (hheeej�%  ]r�%  (jr  ]r�%  (jt  ]r�%  (jv  ]r�%  (hh"e]r�%  (hh	e]r�%  (hjN  e]r�%  (j{  ]r�%  (hhe]r�%  (hh	e]r�%  (hhe]r�%  (j�  ]r�%  (hh	e]r�%  (hh	eeee]r�%  (hheeej�%  j�%  j�%  j�%  j�%  j�%  ]r�%  (jr  ]r�%  (jt  ]r�%  (jv  ]r�%  (hh"e]r�%  (hh	e]r�%  (hjN  e]r�%  (j{  ]r�%  (hhe]r�%  (hh	e]r�%  (hhe]r�%  (j�  ]r�%  (hh	e]r &  (hh	eeee]r&  (hheeej�%  j�%  j�%  j�%  ]r&  (jr  ]r&  (jt  ]r&  (jv  ]r&  (hh"e]r&  (hh	e]r&  (hjN  e]r&  (j{  ]r	&  (hhe]r
&  (hh	e]r&  (hhe]r&  (j�  ]r&  (hh	e]r&  (hh	eeee]r&  (hheee]r&  (jr  ]r&  (jt  ]r&  (jv  ]r&  (hh"e]r&  (hh	e]r&  (hjN  e]r&  (j{  ]r&  (hhe]r&  (hh	e]r&  (hhe]r&  (j�  ]r&  (hh	e]r&  (hh	eeee]r&  (hheee]r&  (jr  ]r&  (jt  ]r &  (jv  ]r!&  (hh"e]r"&  (hh	e]r#&  (hjN  e]r$&  (j{  ]r%&  (hhe]r&&  (hh	e]r'&  (hhe]r(&  (j�  ]r)&  (hh	e]r*&  (hh	eeee]r+&  (hheeej&  j&  j&  j&  j&  j&  j&  j&  j&  j&  j&  j&  ]r,&  (jr  ]r-&  (jt  ]r.&  (jv  ]r/&  (hh"e]r0&  (hh	e]r1&  (hjN  e]r2&  (j{  ]r3&  (hhe]r4&  (hh	e]r5&  (hhe]r6&  (j�  ]r7&  (hh	e]r8&  (hh	eeee]r9&  (hheeej,&  j,&  j,&  j,&  ]r:&  (jr  ]r;&  (jt  ]r<&  (jv  ]r=&  (hh"e]r>&  (hh	e]r?&  (hjN  e]r@&  (j{  ]rA&  (hhe]rB&  (hh	e]rC&  (hhe]rD&  (j�  ]rE&  (hh	e]rF&  (hh	eeee]rG&  (hheeej:&  j:&  ]rH&  (jr  ]rI&  (jt  ]rJ&  (jv  ]rK&  (hh"e]rL&  (hh	e]rM&  (hjN  e]rN&  (j{  ]rO&  (hhe]rP&  (hh	e]rQ&  (hhe]rR&  (j�  ]rS&  (hh	e]rT&  (hh	eeee]rU&  (hheeejH&  jH&  jH&  jH&  jH&  jH&  jH&  ]rV&  (jr  ]rW&  (jt  ]rX&  (jv  ]rY&  (hh"e]rZ&  (hhe]r[&  (hjN  e]r\&  (j{  ]r]&  (hhe]r^&  (hh	e]r_&  (hhe]r`&  (j�  ]ra&  (hh	e]rb&  (hh	eeee]rc&  (hheeejV&  jV&  jV&  ]rd&  (jr  ]re&  (jt  ]rf&  (jv  ]rg&  (hh"e]rh&  (hhe]ri&  (hjN  e]rj&  (j{  ]rk&  (hhe]rl&  (hh	e]rm&  (hhe]rn&  (j�  ]ro&  (hh	e]rp&  (hh	eeee]rq&  (hheee]rr&  (jr  ]rs&  (jt  ]rt&  (jv  ]ru&  (hh"e]rv&  (hhe]rw&  (hjN  e]rx&  (j{  ]ry&  (hhe]rz&  (hh	e]r{&  (hhe]r|&  (j�  ]r}&  (hh	e]r~&  (hh	eeee]r&  (hheeejr&  jr&  jr&  ]r�&  (jr  ]r�&  (jt  ]r�&  (jv  ]r�&  (hh"e]r�&  (hhe]r�&  (hjN  e]r�&  (j{  ]r�&  (hhe]r�&  (hh	e]r�&  (hhe]r�&  (j�  ]r�&  (hh	e]r�&  (hh	eeee]r�&  (hheeej�&  j�&  j�&  ]r�&  (jr  ]r�&  (jt  ]r�&  (jv  ]r�&  (hh"e]r�&  (hhe]r�&  (hjN  e]r�&  (j{  ]r�&  (hhe]r�&  (hh	e]r�&  (hhe]r�&  (j�  ]r�&  (hh	e]r�&  (hh	eeee]r�&  (hheeej�&  j�&  j�&  j�&  j�&  j�&  j�&  j�&  j�&  ]r�&  (jr  ]r�&  (jt  ]r�&  (jv  ]r�&  (hh"e]r�&  (hhe]r�&  (hjN  e]r�&  (j{  ]r�&  (hhe]r�&  (hh	e]r�&  (hhe]r�&  (j�  ]r�&  (hh	e]r�&  (hh	eeee]r�&  (hheeej�&  j�&  j�&  ]r�&  (jr  ]r�&  (jt  ]r�&  (jv  ]r�&  (hh"e]r�&  (hhe]r�&  (hjN  e]r�&  (j{  ]r�&  (hhe]r�&  (hh	e]r�&  (hhe]r�&  (j�  ]r�&  (hh	e]r�&  (hh	eeee]r�&  (hheeej�&  j�&  j�&  j�&  j�&  j�&  ]r�&  (jr  ]r�&  (jt  ]r�&  (jv  ]r�&  (hh"e]r�&  (hhe]r�&  (hjN  e]r�&  (j{  ]r�&  (hhe]r�&  (hh	e]r�&  (hhe]r�&  (j�  ]r�&  (hh	e]r�&  (hh	eeee]r�&  (hheeej�&  j�&  ]r�&  (jr  ]r�&  (jt  ]r�&  (jv  ]r�&  (hh"e]r�&  (hhe]r�&  (hjN  e]r�&  (j{  ]r�&  (hhe]r�&  (hh	e]r�&  (hhe]r�&  (j�  ]r�&  (hh	e]r�&  (hh	eeee]r�&  (hheeej�&  ]r�&  (jr  ]r�&  (jt  ]r�&  (jv  ]r�&  (hh"e]r�&  (hhe]r�&  (hjN  e]r�&  (j{  ]r�&  (hhe]r�&  (hh	e]r�&  (hhe]r�&  (j�  ]r�&  (hh	e]r�&  (hh	eeee]r�&  (hheeej�&  j�&  j�&  j�&  j�&  j�&  j�&  j�&  j�&  ]r�&  (jr  ]r�&  (jt  ]r�&  (jv  ]r�&  (hh"e]r�&  (hhe]r�&  (hjN  e]r�&  (j{  ]r�&  (hhe]r�&  (hh	e]r�&  (hhe]r�&  (j�  ]r�&  (hh	e]r�&  (hh	eeee]r�&  (hheeej�&  ]r�&  (jr  ]r�&  (jt  ]r�&  (jv  ]r�&  (hh"e]r�&  (hhe]r�&  (hjN  e]r�&  (j{  ]r�&  (hhe]r�&  (hh	e]r�&  (hhe]r�&  (j�  ]r�&  (hh	e]r�&  (hh	eeee]r�&  (hheee]r�&  (jr  ]r�&  (jt  ]r '  (jv  ]r'  (hh"e]r'  (hhe]r'  (hjN  e]r'  (j{  ]r'  (hhe]r'  (hh	e]r'  (hhe]r'  (j�  ]r	'  (hh	e]r
'  (hh	eeee]r'  (hheeej�&  ]r'  (jr  ]r'  (jt  ]r'  (jv  ]r'  (hh	e]r'  (hhe]r'  (hjN  e]r'  (j{  ]r'  (hhe]r'  (hh	e]r'  (hhe]r'  (j�  ]r'  (hh	e]r'  (hh	eeee]r'  (hheeej'  j'  j'  j'  j'  ]r'  (jr  ]r'  (jt  ]r'  (jv  ]r'  (hh	e]r'  (hhe]r'  (hjN  e]r '  (j{  ]r!'  (hhe]r"'  (hh	e]r#'  (hhe]r$'  (j�  ]r%'  (hh	e]r&'  (hh	eeee]r''  (hheeej'  j'  ]r('  (jr  ]r)'  (jt  ]r*'  (jv  ]r+'  (hh	e]r,'  (hhe]r-'  (hjN  e]r.'  (j{  ]r/'  (hhe]r0'  (hh	e]r1'  (hhe]r2'  (j�  ]r3'  (hh	e]r4'  (hh	eeee]r5'  (hheeej('  j('  j('  j('  ]r6'  (jr  ]r7'  (jt  ]r8'  (jv  ]r9'  (hh	e]r:'  (hhe]r;'  (hjN  e]r<'  (j{  ]r='  (hhe]r>'  (hh	e]r?'  (hhe]r@'  (j�  ]rA'  (hh	e]rB'  (hh	eeee]rC'  (hheee]rD'  (jr  ]rE'  (jt  ]rF'  (jv  ]rG'  (hh	e]rH'  (hhe]rI'  (hjN  e]rJ'  (j{  ]rK'  (hhe]rL'  (hh	e]rM'  (hhe]rN'  (j�  ]rO'  (hh	e]rP'  (hh	eeee]rQ'  (hheeejD'  jD'  jD'  ]rR'  (jr  ]rS'  (jt  ]rT'  (jv  ]rU'  (hh	e]rV'  (hhe]rW'  (hjN  e]rX'  (j{  ]rY'  (hhe]rZ'  (hh	e]r['  (hhe]r\'  (j�  ]r]'  (hh	e]r^'  (hh	eeee]r_'  (hheeejR'  ]r`'  (jr  ]ra'  (jt  ]rb'  (jv  ]rc'  (hh	e]rd'  (hhe]re'  (hjN  e]rf'  (j{  ]rg'  (hhe]rh'  (hh	e]ri'  (hhe]rj'  (j�  ]rk'  (hh	e]rl'  (hh	eeee]rm'  (hheeej`'  ]rn'  (jr  ]ro'  (jt  ]rp'  (jv  ]rq'  (hh"e]rr'  (hhe]rs'  (hjN  e]rt'  (j{  ]ru'  (hhe]rv'  (hh	e]rw'  (hhe]rx'  (j�  ]ry'  (hh	e]rz'  (hh	eeee]r{'  (hheeejn'  jn'  jn'  jn'  jn'  jn'  jn'  jn'  jn'  jn'  jn'  ]r|'  (jr  ]r}'  (jt  ]r~'  (jv  ]r'  (hh	e]r�'  (hhe]r�'  (hjN  e]r�'  (j{  ]r�'  (hhe]r�'  (hh	e]r�'  (hhe]r�'  (j�  ]r�'  (hh	e]r�'  (hh	eeee]r�'  (hheeej|'  j|'  j|'  ]r�'  (jr  ]r�'  (jt  ]r�'  (jv  ]r�'  (hh	e]r�'  (hhe]r�'  (hjN  e]r�'  (j{  ]r�'  (hhe]r�'  (hh	e]r�'  (hhe]r�'  (j�  ]r�'  (hh	e]r�'  (hh	eeee]r�'  (hheeej�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  ]r�'  (jr  ]r�'  (jt  ]r�'  (jv  ]r�'  (hh	e]r�'  (hhe]r�'  (hjN  e]r�'  (j{  ]r�'  (hhe]r�'  (hh	e]r�'  (hhe]r�'  (j�  ]r�'  (hh	e]r�'  (hh	eeee]r�'  (hheeej�'  j�'  j�'  ]r�'  (jr  ]r�'  (jt  ]r�'  (jv  ]r�'  (hh	e]r�'  (hhe]r�'  (hjN  e]r�'  (j{  ]r�'  (hhe]r�'  (hh	e]r�'  (hhe]r�'  (j�  ]r�'  (hh	e]r�'  (hh	eeee]r�'  (hheeej�'  j�'  j�'  j�'  j�'  ]r�'  (jr  ]r�'  (jt  ]r�'  (jv  ]r�'  (hh	e]r�'  (hhe]r�'  (hjN  e]r�'  (j{  ]r�'  (hhe]r�'  (hh	e]r�'  (hhe]r�'  (j�  ]r�'  (hh	e]r�'  (hh	eeee]r�'  (hheeej�'  ]r�'  (jr  ]r�'  (jt  ]r�'  (jv  ]r�'  (hh	e]r�'  (hhe]r�'  (hjN  e]r�'  (j{  ]r�'  (hhe]r�'  (hh	e]r�'  (hhe]r�'  (j�  ]r�'  (hh	e]r�'  (hh	eeee]r�'  (hheeej�'  j�'  j�'  ]r�'  (jr  ]r�'  (jt  ]r�'  (jv  ]r�'  (hh	e]r�'  (hhe]r�'  (hjN  e]r�'  (j{  ]r�'  (hhe]r�'  (hh	e]r�'  (hhe]r�'  (j�  ]r�'  (hh	e]r�'  (hh	eeee]r�'  (hheeej�'  ]r�'  (jr  ]r�'  (jt  ]r�'  (jv  ]r�'  (hh"e]r�'  (hhe]r�'  (hjN  e]r�'  (j{  ]r�'  (hhe]r�'  (hh	e]r�'  (hhe]r�'  (j�  ]r�'  (hh	e]r�'  (hh	eeee]r�'  (hheeej�'  j�'  j�'  j�'  j�'  j�'  ]r�'  (jr  ]r�'  (jt  ]r�'  (jv  ]r�'  (hh"e]r�'  (hh	e]r�'  (hjN  e]r�'  (j{  ]r�'  (hhe]r�'  (hh	e]r�'  (hhe]r�'  (j�  ]r�'  (hh	e]r�'  (hh	eeee]r�'  (hheeej�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  ]r�'  (jr  ]r�'  (jt  ]r�'  (jv  ]r�'  (hh"e]r�'  (hh	e]r�'  (hjN  e]r (  (j{  ]r(  (hhe]r(  (hh	e]r(  (hhe]r(  (j�  ]r(  (hh	e]r(  (hh	eeee]r(  (hheeej�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  ]r(  (jr  ]r	(  (jt  ]r
(  (jv  ]r(  (hh"e]r(  (hh	e]r(  (hjN  e]r(  (j{  ]r(  (hhe]r(  (hh	e]r(  (hhe]r(  (j�  ]r(  (hh	e]r(  (hh	eeee]r(  (hheeej(  j(  ]r(  (jr  ]r(  (jt  ]r(  (jv  ]r(  (hh"e]r(  (hh	e]r(  (hjN  e]r(  (j{  ]r(  (hhe]r(  (hh	e]r(  (hhe]r (  (j�  ]r!(  (hh	e]r"(  (hh	eeee]r#(  (hheeej(  j(  j(  ]r$(  (jr  ]r%(  (jt  ]r&(  (jv  ]r'(  (hh"e]r((  (hh	e]r)(  (hjN  e]r*(  (j{  ]r+(  (hhe]r,(  (hh	e]r-(  (hhe]r.(  (j�  ]r/(  (hh	e]r0(  (hh	eeee]r1(  (hheeej$(  j$(  j$(  j$(  j$(  ]r2(  (jr  ]r3(  (jt  ]r4(  (jv  ]r5(  (hh"e]r6(  (hh	e]r7(  (hjN  e]r8(  (j{  ]r9(  (hhe]r:(  (hh	e]r;(  (hhe]r<(  (j�  ]r=(  (hh	e]r>(  (hh	eeee]r?(  (hheeej2(  j2(  j2(  j2(  j2(  j2(  j2(  j2(  j2(  ]r@(  (jr  ]rA(  (jt  ]rB(  (jv  ]rC(  (hh"e]rD(  (hh	e]rE(  (hjN  e]rF(  (j{  ]rG(  (hhe]rH(  (hh	e]rI(  (hhe]rJ(  (j�  ]rK(  (hh	e]rL(  (hh	eeee]rM(  (hheeej@(  j@(  ]rN(  (jr  ]rO(  (jt  ]rP(  (jv  ]rQ(  (hh"e]rR(  (hh	e]rS(  (hjN  e]rT(  (j{  ]rU(  (hhe]rV(  (hh	e]rW(  (hhe]rX(  (j�  ]rY(  (hh	e]rZ(  (hh	eeee]r[(  (hheeejN(  ]r\(  (jr  ]r](  (jt  ]r^(  (jv  ]r_(  (hh"e]r`(  (hh	e]ra(  (hjN  e]rb(  (j{  ]rc(  (hhe]rd(  (hh	e]re(  (hhe]rf(  (j�  ]rg(  (hh	e]rh(  (hh	eeee]ri(  (hheeej\(  j\(  j\(  ]rj(  (jr  ]rk(  (jt  ]rl(  (jv  ]rm(  (hh"e]rn(  (hh	e]ro(  (hjN  e]rp(  (j{  ]rq(  (hhe]rr(  (hh	e]rs(  (hhe]rt(  (j�  ]ru(  (hh	e]rv(  (hh	eeee]rw(  (hheeejj(  jj(  ]rx(  (jr  ]ry(  (jt  ]rz(  (jv  ]r{(  (hh"e]r|(  (hh	e]r}(  (hjN  e]r~(  (j{  ]r(  (hhe]r�(  (hh	e]r�(  (hhe]r�(  (j�  ]r�(  (hh	e]r�(  (hh	eeee]r�(  (hheeejx(  jx(  ]r�(  (jr  ]r�(  (jt  ]r�(  (jv  ]r�(  (hh"e]r�(  (hh	e]r�(  (hjN  e]r�(  (j{  ]r�(  (hhe]r�(  (hh	e]r�(  (hhe]r�(  (j�  ]r�(  (hh	e]r�(  (hh	eeee]r�(  (hheeej�(  j�(  j�(  j�(  j�(  j�(  j�(  ]r�(  (jr  ]r�(  (jt  ]r�(  (jv  ]r�(  (hh"e]r�(  (hh	e]r�(  (hjN  e]r�(  (j{  ]r�(  (hhe]r�(  (hh	e]r�(  (hhe]r�(  (j�  ]r�(  (hh	e]r�(  (hh	eeee]r�(  (hheeej�(  j�(  j�(  j�(  ]r�(  (jr  ]r�(  (jt  ]r�(  (jv  ]r�(  (hh"e]r�(  (hh	e]r�(  (hjN  e]r�(  (j{  ]r�(  (hhe]r�(  (hh	e]r�(  (hhe]r�(  (j�  ]r�(  (hh	e]r�(  (hh	eeee]r�(  (hheeej�(  ]r�(  (jr  ]r�(  (jt  ]r�(  (jv  ]r�(  (hh"e]r�(  (hh	e]r�(  (hjN  e]r�(  (j{  ]r�(  (hhe]r�(  (hh	e]r�(  (hhe]r�(  (j�  ]r�(  (hh	e]r�(  (hh	eeee]r�(  (hheeej�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  ]r�(  (jr  ]r�(  (jt  ]r�(  (jv  ]r�(  (hh"e]r�(  (hh	e]r�(  (hjN  e]r�(  (j{  ]r�(  (hhe]r�(  (hh	e]r�(  (hhe]r�(  (j�  ]r�(  (hh	e]r�(  (hh	eeee]r�(  (hheeej�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  ]r�(  (jr  ]r�(  (jt  ]r�(  (jv  ]r�(  (hh"e]r�(  (hh	e]r�(  (hjN  e]r�(  (j{  ]r�(  (hhe]r�(  (hh	e]r�(  (hhe]r�(  (j�  ]r�(  (hh	e]r�(  (hh	eeee]r�(  (hheeej�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  ]r�(  (jr  ]r�(  (jt  ]r�(  (jv  ]r�(  (hh"e]r�(  (hh	e]r�(  (hjN  e]r�(  (j{  ]r�(  (hhe]r�(  (hh	e]r�(  (hhe]r�(  (j�  ]r�(  (hh	e]r�(  (hh	eeee]r�(  (hheeej�(  j�(  ]r�(  (jr  ]r�(  (jt  ]r�(  (jv  ]r�(  (hh"e]r�(  (hh	e]r�(  (hjN  e]r�(  (j{  ]r�(  (hhe]r�(  (hh	e]r�(  (hhe]r�(  (j�  ]r�(  (hh	e]r�(  (hh	eeee]r�(  (hheeej�(  ]r�(  (jr  ]r�(  (jt  ]r�(  (jv  ]r�(  (hh"e]r�(  (hh	e]r�(  (hjN  e]r�(  (j{  ]r�(  (hhe]r�(  (hh	e]r�(  (hhe]r )  (j�  ]r)  (hh	e]r)  (hh	eeee]r)  (hheeej�(  j�(  j�(  j�(  j�(  j�(  ]r)  (jr  ]r)  (jt  ]r)  (jv  ]r)  (hh"e]r)  (hh	e]r	)  (hjN  e]r
)  (j{  ]r)  (hhe]r)  (hh	e]r)  (hhe]r)  (j�  ]r)  (hh	e]r)  (hh	eeee]r)  (hheeej)  ]r)  (jr  ]r)  (jt  ]r)  (jv  ]r)  (hh"e]r)  (hh	e]r)  (hjN  e]r)  (j{  ]r)  (hhe]r)  (hh	e]r)  (hhe]r)  (j�  ]r)  (hh	e]r)  (hh	eeee]r)  (hheeej)  j)  j)  j)  j)  j)  j)  j)  ]r )  (jr  ]r!)  (jt  ]r")  (jv  ]r#)  (hh"e]r$)  (hh	e]r%)  (hjN  e]r&)  (j{  ]r')  (hhe]r()  (hh	e]r))  (hhe]r*)  (j�  ]r+)  (hh	e]r,)  (hh	eeee]r-)  (hheee]r.)  (jr  ]r/)  (jt  ]r0)  (jv  ]r1)  (hh"e]r2)  (hh	e]r3)  (hjN  e]r4)  (j{  ]r5)  (hhe]r6)  (hh	e]r7)  (hhe]r8)  (j�  ]r9)  (hh	e]r:)  (hh	eeee]r;)  (hheeej.)  j.)  j.)  j.)  j.)  j.)  ]r<)  (jr  ]r=)  (jt  ]r>)  (jv  ]r?)  (hh"e]r@)  (hh	e]rA)  (hjN  e]rB)  (j{  ]rC)  (hhe]rD)  (hh	e]rE)  (hhe]rF)  (j�  ]rG)  (hh	e]rH)  (hh	eeee]rI)  (hheeej<)  j<)  j<)  j<)  j<)  j<)  j<)  j<)  j<)  ]rJ)  (jr  ]rK)  (jt  ]rL)  (jv  ]rM)  (hh"e]rN)  (hh	e]rO)  (hjN  e]rP)  (j{  ]rQ)  (hhe]rR)  (hh	e]rS)  (hhe]rT)  (j�  ]rU)  (hh	e]rV)  (hh	eeee]rW)  (hheeejJ)  jJ)  jJ)  ]rX)  (jr  ]rY)  (jt  ]rZ)  (jv  ]r[)  (hh"e]r\)  (hh	e]r])  (hjN  e]r^)  (j{  ]r_)  (hhe]r`)  (hh	e]ra)  (hhe]rb)  (j�  ]rc)  (hh	e]rd)  (hh	eeee]re)  (hheeejX)  jX)  jX)  jX)  ]rf)  (jr  ]rg)  (jt  ]rh)  (jv  ]ri)  (hh"e]rj)  (hh	e]rk)  (hjN  e]rl)  (j{  ]rm)  (hhe]rn)  (hh	e]ro)  (hhe]rp)  (j�  ]rq)  (hh	e]rr)  (hh	eeee]rs)  (hheeejf)  jf)  jf)  ]rt)  (jr  ]ru)  (jt  ]rv)  (jv  ]rw)  (hh"e]rx)  (hh	e]ry)  (hjN  e]rz)  (j{  ]r{)  (hhe]r|)  (hh	e]r})  (hhe]r~)  (j�  ]r)  (hh	e]r�)  (hh	eeee]r�)  (hheeejt)  jt)  jt)  jt)  jt)  jt)  jt)  jt)  jt)  jt)  ]r�)  (jr  ]r�)  (jt  ]r�)  (jv  ]r�)  (hh"e]r�)  (hh	e]r�)  (hjN  e]r�)  (j{  ]r�)  (hhe]r�)  (hh	e]r�)  (hhe]r�)  (j�  ]r�)  (hh	e]r�)  (hh	eeee]r�)  (hheeej�)  j�)  j�)  ]r�)  (jr  ]r�)  (jt  ]r�)  (jv  ]r�)  (hh"e]r�)  (hh	e]r�)  (hjN  e]r�)  (j{  ]r�)  (hhe]r�)  (hh	e]r�)  (hhe]r�)  (j�  ]r�)  (hh	e]r�)  (hh	eeee]r�)  (hheee]r�)  (jr  ]r�)  (jt  ]r�)  (jv  ]r�)  (hh"e]r�)  (hh	e]r�)  (hjN  e]r�)  (j{  ]r�)  (hhe]r�)  (hh	e]r�)  (hhe]r�)  (j�  ]r�)  (hh	e]r�)  (hh	eeee]r�)  (hheeej�)  j�)  ]r�)  (jr  ]r�)  (jt  ]r�)  (jv  ]r�)  (hh"e]r�)  (hh	e]r�)  (hjN  e]r�)  (j{  ]r�)  (hhe]r�)  (hh	e]r�)  (hhe]r�)  (j�  ]r�)  (hh	e]r�)  (hh	eeee]r�)  (hheeej�)  j�)  j�)  ]r�)  (jr  ]r�)  (jt  ]r�)  (jv  ]r�)  (hh"e]r�)  (hhe]r�)  (hjN  e]r�)  (j{  ]r�)  (hhe]r�)  (hh	e]r�)  (hhe]r�)  (j�  ]r�)  (hh	e]r�)  (hh	eeee]r�)  (hheeej�)  j�)  j�)  j�)  j�)  j�)  j�)  ]r�)  (jr  ]r�)  (X   Oblr�)  ]r�)  (j^  ]r�)  (hh	e]r�)  (hhe]r�)  (hh&e]r�)  (j^  ]r�)  (hX   rr�)  e]r�)  (hX   circler�)  e]r�)  (hh&e]r�)  (X	   Next-Mover�)  ]r�)  (hhe]r�)  (hheeee]r�)  (hh&eee]r�)  (jr  ]r�)  (j�)  ]r�)  (j^  ]r�)  (hh	e]r�)  (hhe]r�)  (hh&e]r�)  (j^  ]r�)  (hj�)  e]r�)  (hj�)  e]r�)  (hh&e]r�)  (j�)  ]r�)  (hhe]r�)  (hheeee]r�)  (hh&eeej�)  j�)  j�)  j�)  ]r�)  (jr  ]r�)  (j�)  ]r�)  (j^  ]r�)  (hh	e]r�)  (hhe]r�)  (hh&e]r�)  (j^  ]r�)  (hj�)  e]r�)  (hh	e]r�)  (hh&e]r�)  (j�)  ]r�)  (hhe]r�)  (hheeee]r�)  (hh&eeej�)  ]r�)  (jr  ]r�)  (j�)  ]r�)  (j^  ]r�)  (hh	e]r�)  (hhe]r�)  (hh&e]r�)  (j^  ]r�)  (hh	e]r�)  (hh	e]r�)  (hh&e]r *  (j�)  ]r*  (hhe]r*  (hheeee]r*  (hh&eeej�)  j�)  j�)  ]r*  (jr  ]r*  (j�)  ]r*  (j^  ]r*  (hh	e]r*  (hhe]r	*  (hh&e]r
*  (j^  ]r*  (hh	e]r*  (hh	e]r*  (hh&e]r*  (j�)  ]r*  (hhe]r*  (hheeee]r*  (hh&eeej*  j*  j*  j*  j*  j*  j*  ]r*  (jr  ]r*  (j�)  ]r*  (j^  ]r*  (hh	e]r*  (hhe]r*  (hh&e]r*  (j^  ]r*  (hh	e]r*  (hh	e]r*  (hh&e]r*  (j�)  ]r*  (hhe]r*  (hheeee]r*  (hh&eee]r *  (jr  ]r!*  (j�)  ]r"*  (j^  ]r#*  (hh	e]r$*  (hhe]r%*  (hh&e]r&*  (j^  ]r'*  (hh	e]r(*  (hh	e]r)*  (hh&e]r**  (j�)  ]r+*  (hhe]r,*  (hheeee]r-*  (hh&eeej *  j *  j *  j *  j *  j *  ]r.*  (jr  ]r/*  (j�)  ]r0*  (j^  ]r1*  (hh	e]r2*  (hhe]r3*  (hh&e]r4*  (j^  ]r5*  (hh	e]r6*  (hh	e]r7*  (hh&e]r8*  (j�)  ]r9*  (hhe]r:*  (hheeee]r;*  (hh&eeej.*  j.*  j.*  j.*  j.*  j.*  j.*  ]r<*  (jr  ]r=*  (j�)  ]r>*  (j^  ]r?*  (hh	e]r@*  (hhe]rA*  (hh&e]rB*  (j^  ]rC*  (hh	e]rD*  (hh	e]rE*  (hh&e]rF*  (j�)  ]rG*  (hhe]rH*  (hheeee]rI*  (hh&eeej<*  ]rJ*  (jr  ]rK*  (j�)  ]rL*  (j^  ]rM*  (hh	e]rN*  (hhe]rO*  (hh&e]rP*  (j^  ]rQ*  (hh	e]rR*  (hh	e]rS*  (hh&e]rT*  (j�)  ]rU*  (hhe]rV*  (hheeee]rW*  (hh&eeejJ*  jJ*  jJ*  jJ*  ]rX*  (jr  ]rY*  (j�)  ]rZ*  (j^  ]r[*  (hh	e]r\*  (hh	e]r]*  (hh&e]r^*  (j^  ]r_*  (hh	e]r`*  (hh	e]ra*  (hh&e]rb*  (j�)  ]rc*  (hhe]rd*  (hheeee]re*  (hh&eeejX*  jX*  ]rf*  (jr  ]rg*  (j�)  ]rh*  (j^  ]ri*  (hh	e]rj*  (hh	e]rk*  (hh&e]rl*  (j^  ]rm*  (hh	e]rn*  (hh	e]ro*  (hh&e]rp*  (j�)  ]rq*  (hhe]rr*  (hheeee]rs*  (hh&eeejf*  jf*  jf*  jf*  jf*  e(]rt*  (X   Normsru*  ]rv*  (X   Oblrw*  ]rx*  (X   Movedry*  ]rz*  (hh	e]r{*  (hh	e]r|*  (hjN  e]r}*  (X   Movedr~*  ]r*  (hh	e]r�*  (hhe]r�*  (hjN  e]r�*  (X	   Next-Mover�*  ]r�*  (hh	e]r�*  (hh	eeee]r�*  (hh&ee]r�*  (h]r�*  (hh e]r�*  (hhe]r�*  (hh	e]r�*  (h%heeejt*  jt*  jt*  jt*  jt*  jt*  jt*  jt*  ]r�*  (ju*  ]r�*  (jw*  ]r�*  (jy*  ]r�*  (hh	e]r�*  (hh	e]r�*  (hjN  e]r�*  (j~*  ]r�*  (hh	e]r�*  (hhe]r�*  (hjN  e]r�*  (j�*  ]r�*  (hh	e]r�*  (hh	eeee]r�*  (hh&ee]r�*  (h]r�*  (hh e]r�*  (hhe]r�*  (hh	e]r�*  (h%heee]r�*  (ju*  ]r�*  (jw*  ]r�*  (jy*  ]r�*  (hh	e]r�*  (hh	e]r�*  (hjN  e]r�*  (j~*  ]r�*  (hh	e]r�*  (hhe]r�*  (hjN  e]r�*  (j�*  ]r�*  (hh	e]r�*  (hh	eeee]r�*  (hh&ee]r�*  (h]r�*  (hh e]r�*  (hhe]r�*  (hh	e]r�*  (h%heeej�*  j�*  j�*  j�*  ]r�*  (ju*  ]r�*  (jw*  ]r�*  (jy*  ]r�*  (hh	e]r�*  (hh	e]r�*  (hjN  e]r�*  (j~*  ]r�*  (hh	e]r�*  (hhe]r�*  (hjN  e]r�*  (j�*  ]r�*  (hh	e]r�*  (hh	eeee]r�*  (hh&ee]r�*  (h]r�*  (hh e]r�*  (hhe]r�*  (hh	e]r�*  (h%heeej�*  j�*  j�*  j�*  j�*  j�*  j�*  ]r�*  (ju*  ]r�*  (jw*  ]r�*  (jy*  ]r�*  (hh	e]r�*  (hh	e]r�*  (hjN  e]r�*  (j~*  ]r�*  (hh	e]r�*  (hhe]r�*  (hjN  e]r�*  (j�*  ]r�*  (hh	e]r�*  (hh	eeee]r�*  (hh&ee]r�*  (h]r�*  (hh e]r�*  (hhe]r�*  (hh	e]r�*  (h%heee]r�*  (ju*  ]r�*  (jw*  ]r�*  (jy*  ]r�*  (hh	e]r�*  (hh	e]r�*  (hjN  e]r�*  (j~*  ]r�*  (hh	e]r�*  (hhe]r�*  (hjN  e]r�*  (j�*  ]r�*  (hh	e]r�*  (hh	eeee]r�*  (hh&ee]r�*  (h]r�*  (hh e]r�*  (hhe]r�*  (hh	e]r�*  (h%heeej�*  j�*  ]r�*  (ju*  ]r�*  (jw*  ]r�*  (jy*  ]r�*  (hh	e]r�*  (hh	e]r�*  (hjN  e]r�*  (j~*  ]r�*  (hh	e]r�*  (hhe]r�*  (hjN  e]r�*  (j�*  ]r�*  (hh	e]r�*  (hh	eeee]r�*  (hh&ee]r�*  (h]r�*  (hh e]r�*  (hhe]r�*  (hh	e]r�*  (h%heee]r�*  (ju*  ]r�*  (jw*  ]r +  (jy*  ]r+  (hh	e]r+  (hh	e]r+  (hjN  e]r+  (j~*  ]r+  (hh	e]r+  (hhe]r+  (hjN  e]r+  (j�*  ]r	+  (hh	e]r
+  (hh	eeee]r+  (hh&ee]r+  (h]r+  (hh e]r+  (hhe]r+  (hh	e]r+  (h%heee]r+  (ju*  ]r+  (jw*  ]r+  (jy*  ]r+  (hh	e]r+  (hh	e]r+  (hjN  e]r+  (j~*  ]r+  (hh	e]r+  (hhe]r+  (hjN  e]r+  (j�*  ]r+  (hh	e]r+  (hh	eeee]r+  (hh&ee]r+  (h]r +  (hh e]r!+  (hhe]r"+  (hh	e]r#+  (h%heeej+  j+  ]r$+  (ju*  ]r%+  (jw*  ]r&+  (jy*  ]r'+  (hh	e]r(+  (hh	e]r)+  (hjN  e]r*+  (j~*  ]r++  (hh	e]r,+  (hhe]r-+  (hjN  e]r.+  (j�*  ]r/+  (hh	e]r0+  (hh	eeee]r1+  (hh&ee]r2+  (h]r3+  (hh e]r4+  (hhe]r5+  (hh	e]r6+  (h%heeej$+  j$+  j$+  j$+  j$+  j$+  j$+  j$+  j$+  j$+  j$+  j$+  ]r7+  (ju*  ]r8+  (jw*  ]r9+  (jy*  ]r:+  (hh	e]r;+  (hh	e]r<+  (hjN  e]r=+  (j~*  ]r>+  (hh	e]r?+  (hhe]r@+  (hjN  e]rA+  (j�*  ]rB+  (hh	e]rC+  (hh	eeee]rD+  (hh&ee]rE+  (h]rF+  (hh e]rG+  (hhe]rH+  (hh	e]rI+  (h%heeej7+  j7+  j7+  j7+  j7+  j7+  j7+  j7+  j7+  ]rJ+  (ju*  ]rK+  (jw*  ]rL+  (jy*  ]rM+  (hh	e]rN+  (hh	e]rO+  (hjN  e]rP+  (j~*  ]rQ+  (hh	e]rR+  (hhe]rS+  (hjN  e]rT+  (j�*  ]rU+  (hh	e]rV+  (hh	eeee]rW+  (hh&ee]rX+  (h]rY+  (hh e]rZ+  (hhe]r[+  (hh	e]r\+  (h%heeejJ+  jJ+  jJ+  jJ+  jJ+  jJ+  ]r]+  (ju*  ]r^+  (jw*  ]r_+  (jy*  ]r`+  (hh	e]ra+  (hh	e]rb+  (hjN  e]rc+  (j~*  ]rd+  (hh	e]re+  (hhe]rf+  (hjN  e]rg+  (j�*  ]rh+  (hh	e]ri+  (hh	eeee]rj+  (hh&ee]rk+  (h]rl+  (hh e]rm+  (hhe]rn+  (hh	e]ro+  (h%heeej]+  ]rp+  (ju*  ]rq+  (jw*  ]rr+  (jy*  ]rs+  (hh	e]rt+  (hh	e]ru+  (hjN  e]rv+  (j~*  ]rw+  (hhe]rx+  (hhe]ry+  (hjN  e]rz+  (j�*  ]r{+  (hh	e]r|+  (hh	eeee]r}+  (hh&ee]r~+  (h]r+  (hh e]r�+  (hhe]r�+  (hh	e]r�+  (h%heeejp+  jp+  jp+  jp+  jp+  jp+  jp+  jp+  jp+  jp+  ]r�+  (ju*  ]r�+  (jw*  ]r�+  (jy*  ]r�+  (hh	e]r�+  (hh	e]r�+  (hjN  e]r�+  (j~*  ]r�+  (hhe]r�+  (hhe]r�+  (hjN  e]r�+  (j�*  ]r�+  (hh	e]r�+  (hh	eeee]r�+  (hh&ee]r�+  (h]r�+  (hh e]r�+  (hhe]r�+  (hh	e]r�+  (h%heeej�+  j�+  ]r�+  (ju*  ]r�+  (jw*  ]r�+  (jy*  ]r�+  (hh	e]r�+  (hh	e]r�+  (hjN  e]r�+  (j~*  ]r�+  (hhe]r�+  (hhe]r�+  (hjN  e]r�+  (j�*  ]r�+  (hh	e]r�+  (hh	eeee]r�+  (hh&ee]r�+  (h]r�+  (hh e]r�+  (hhe]r�+  (hhe]r�+  (h%heee]r�+  (ju*  ]r�+  (jw*  ]r�+  (jy*  ]r�+  (hh	e]r�+  (hh	e]r�+  (hjN  e]r�+  (j~*  ]r�+  (hhe]r�+  (hhe]r�+  (hjN  e]r�+  (j�*  ]r�+  (hh	e]r�+  (hh	eeee]r�+  (hh&ee]r�+  (h]r�+  (hh e]r�+  (hhe]r�+  (hhe]r�+  (h%heeej�+  ]r�+  (ju*  ]r�+  (jw*  ]r�+  (jy*  ]r�+  (hh	e]r�+  (hh	e]r�+  (hjN  e]r�+  (j~*  ]r�+  (hhe]r�+  (hhe]r�+  (hjN  e]r�+  (j�*  ]r�+  (hh	e]r�+  (hh	eeee]r�+  (hh&ee]r�+  (h]r�+  (hh e]r�+  (hhe]r�+  (hhe]r�+  (h%heeej�+  j�+  j�+  j�+  j�+  ]r�+  (ju*  ]r�+  (jw*  ]r�+  (jy*  ]r�+  (hh	e]r�+  (hh	e]r�+  (hjN  e]r�+  (j~*  ]r�+  (hhe]r�+  (hhe]r�+  (hjN  e]r�+  (j�*  ]r�+  (hh	e]r�+  (hh	eeee]r�+  (hh&ee]r�+  (h]r�+  (hh e]r�+  (hhe]r�+  (hhe]r�+  (h%heeej�+  j�+  ]r�+  (ju*  ]r�+  (jw*  ]r�+  (jy*  ]r�+  (hh	e]r�+  (hh	e]r�+  (hjN  e]r�+  (j~*  ]r�+  (hhe]r�+  (hhe]r�+  (hjN  e]r�+  (j�*  ]r�+  (hh	e]r�+  (hh	eeee]r�+  (hh&ee]r�+  (h]r�+  (hh e]r�+  (hhe]r�+  (hhe]r�+  (h%heeej�+  ]r�+  (ju*  ]r�+  (jw*  ]r�+  (jy*  ]r�+  (hh	e]r�+  (hh	e]r�+  (hjN  e]r�+  (j~*  ]r�+  (hhe]r�+  (hhe]r�+  (hjN  e]r�+  (j�*  ]r ,  (hh	e]r,  (hh	eeee]r,  (hh&ee]r,  (h]r,  (hh e]r,  (hhe]r,  (hh	e]r,  (h%heee]r,  (ju*  ]r	,  (jw*  ]r
,  (jy*  ]r,  (hh	e]r,  (hh	e]r,  (hjN  e]r,  (j~*  ]r,  (hhe]r,  (hhe]r,  (hjN  e]r,  (j�*  ]r,  (hh	e]r,  (hh	eeee]r,  (hh&ee]r,  (h]r,  (hh e]r,  (hhe]r,  (hh	e]r,  (h%heeej,  j,  ]r,  (ju*  ]r,  (jw*  ]r,  (jy*  ]r,  (hh	e]r,  (hh	e]r ,  (hjN  e]r!,  (j~*  ]r",  (hhe]r#,  (hhe]r$,  (hjN  e]r%,  (j�*  ]r&,  (hh	e]r',  (hh	eeee]r(,  (hh&ee]r),  (h]r*,  (hh e]r+,  (hhe]r,,  (hh	e]r-,  (h%heeej,  j,  j,  j,  j,  j,  j,  j,  j,  j,  j,  j,  j,  j,  j,  j,  j,  ]r.,  (ju*  ]r/,  (jw*  ]r0,  (jy*  ]r1,  (hh	e]r2,  (hh	e]r3,  (hjN  e]r4,  (j~*  ]r5,  (hhe]r6,  (hhe]r7,  (hjN  e]r8,  (j�*  ]r9,  (hh	e]r:,  (hh	eeee]r;,  (hh&ee]r<,  (h]r=,  (hh e]r>,  (hhe]r?,  (hh	e]r@,  (h%heee]rA,  (ju*  ]rB,  (jw*  ]rC,  (jy*  ]rD,  (hh	e]rE,  (hh	e]rF,  (hjN  e]rG,  (j~*  ]rH,  (hhe]rI,  (hhe]rJ,  (hjN  e]rK,  (j�*  ]rL,  (hh	e]rM,  (hh	eeee]rN,  (hh&ee]rO,  (h]rP,  (hh e]rQ,  (hhe]rR,  (hh	e]rS,  (h%heeejA,  ]rT,  (ju*  ]rU,  (jw*  ]rV,  (jy*  ]rW,  (hh	e]rX,  (hh	e]rY,  (hjN  e]rZ,  (j~*  ]r[,  (hhe]r\,  (hhe]r],  (hjN  e]r^,  (j�*  ]r_,  (hh	e]r`,  (hh	eeee]ra,  (hh&ee]rb,  (h]rc,  (hh e]rd,  (hhe]re,  (hh	e]rf,  (h%heee]rg,  (ju*  ]rh,  (jw*  ]ri,  (jy*  ]rj,  (hh	e]rk,  (hh	e]rl,  (hjN  e]rm,  (j~*  ]rn,  (hhe]ro,  (hhe]rp,  (hjN  e]rq,  (j�*  ]rr,  (hh	e]rs,  (hh	eeee]rt,  (hh&ee]ru,  (h]rv,  (hh e]rw,  (hhe]rx,  (hh	e]ry,  (h%heeejg,  jg,  jg,  ]rz,  (ju*  ]r{,  (jw*  ]r|,  (jy*  ]r},  (hh	e]r~,  (hh	e]r,  (hjN  e]r�,  (j~*  ]r�,  (hhe]r�,  (hhe]r�,  (hjN  e]r�,  (j�*  ]r�,  (hh	e]r�,  (hh	eeee]r�,  (hh&ee]r�,  (h]r�,  (hh e]r�,  (hhe]r�,  (hhe]r�,  (h%heeejz,  jz,  jz,  ]r�,  (ju*  ]r�,  (jw*  ]r�,  (jy*  ]r�,  (hh	e]r�,  (hh	e]r�,  (hjN  e]r�,  (j~*  ]r�,  (hhe]r�,  (hhe]r�,  (hjN  e]r�,  (j�*  ]r�,  (hh	e]r�,  (hh	eeee]r�,  (hh&ee]r�,  (h]r�,  (hh e]r�,  (hhe]r�,  (hhe]r�,  (h%heeej�,  ]r�,  (ju*  ]r�,  (jw*  ]r�,  (jy*  ]r�,  (hh	e]r�,  (hh	e]r�,  (hjN  e]r�,  (j~*  ]r�,  (hhe]r�,  (hhe]r�,  (hjN  e]r�,  (j�*  ]r�,  (hh	e]r�,  (hh	eeee]r�,  (hh&ee]r�,  (h]r�,  (hh e]r�,  (hhe]r�,  (hhe]r�,  (h%heeej�,  ]r�,  (ju*  ]r�,  (jw*  ]r�,  (jy*  ]r�,  (hh	e]r�,  (hh	e]r�,  (hjN  e]r�,  (j~*  ]r�,  (hhe]r�,  (hhe]r�,  (hjN  e]r�,  (j�*  ]r�,  (hh	e]r�,  (hh	eeee]r�,  (hh&ee]r�,  (h]r�,  (hh e]r�,  (hhe]r�,  (hhe]r�,  (h%heeej�,  j�,  j�,  ]r�,  (ju*  ]r�,  (jw*  ]r�,  (jy*  ]r�,  (hh	e]r�,  (hh	e]r�,  (hjN  e]r�,  (j~*  ]r�,  (hhe]r�,  (hhe]r�,  (hjN  e]r�,  (j�*  ]r�,  (hh	e]r�,  (hh	eeee]r�,  (hh&ee]r�,  (h]r�,  (hh e]r�,  (hhe]r�,  (hhe]r�,  (h%heeej�,  j�,  ]r�,  (ju*  ]r�,  (jw*  ]r�,  (jy*  ]r�,  (hh	e]r�,  (hh	e]r�,  (hjN  e]r�,  (j~*  ]r�,  (hhe]r�,  (hhe]r�,  (hjN  e]r�,  (j�*  ]r�,  (hh	e]r�,  (hh	eeee]r�,  (hh&ee]r�,  (h]r�,  (hh e]r�,  (hhe]r�,  (hhe]r�,  (h%heeej�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  ]r�,  (ju*  ]r�,  (jw*  ]r�,  (jy*  ]r�,  (hh	e]r�,  (hh	e]r�,  (hjN  e]r�,  (j~*  ]r�,  (hhe]r�,  (hhe]r�,  (hjN  e]r�,  (j�*  ]r�,  (hh	e]r�,  (hh	eeee]r�,  (hh&ee]r�,  (h]r�,  (hh e]r�,  (hhe]r�,  (hhe]r�,  (h%heee]r�,  (ju*  ]r -  (jw*  ]r-  (jy*  ]r-  (hh	e]r-  (hh	e]r-  (hjN  e]r-  (j~*  ]r-  (hhe]r-  (hhe]r-  (hjN  e]r	-  (j�*  ]r
-  (hh	e]r-  (hh	eeee]r-  (hh&ee]r-  (h]r-  (hh e]r-  (hhe]r-  (hhe]r-  (h%heee]r-  (ju*  ]r-  (jw*  ]r-  (jy*  ]r-  (hh	e]r-  (hh	e]r-  (hjN  e]r-  (j~*  ]r-  (hhe]r-  (hhe]r-  (hjN  e]r-  (j�*  ]r-  (hh	e]r-  (hh	eeee]r-  (hh&ee]r -  (h]r!-  (hh e]r"-  (hhe]r#-  (hhe]r$-  (h%heeej-  j-  ]r%-  (ju*  ]r&-  (jw*  ]r'-  (jy*  ]r(-  (hh	e]r)-  (hh	e]r*-  (hjN  e]r+-  (j~*  ]r,-  (hhe]r--  (hhe]r.-  (hjN  e]r/-  (j�*  ]r0-  (hh	e]r1-  (hh	eeee]r2-  (hh&ee]r3-  (h]r4-  (hh e]r5-  (hhe]r6-  (hhe]r7-  (h%heeej%-  j%-  j%-  j%-  j%-  j%-  j%-  j%-  j%-  ]r8-  (ju*  ]r9-  (jw*  ]r:-  (jy*  ]r;-  (hh	e]r<-  (hh	e]r=-  (hjN  e]r>-  (j~*  ]r?-  (hhe]r@-  (hhe]rA-  (hjN  e]rB-  (j�*  ]rC-  (hh	e]rD-  (hh	eeee]rE-  (hh&ee]rF-  (h]rG-  (hh e]rH-  (hhe]rI-  (hhe]rJ-  (h%heeej8-  j8-  j8-  j8-  ]rK-  (ju*  ]rL-  (jw*  ]rM-  (jy*  ]rN-  (hh	e]rO-  (hh	e]rP-  (hjN  e]rQ-  (j~*  ]rR-  (hhe]rS-  (hhe]rT-  (hjN  e]rU-  (j�*  ]rV-  (hh	e]rW-  (hh	eeee]rX-  (hh&ee]rY-  (h]rZ-  (hh e]r[-  (hhe]r\-  (hhe]r]-  (h%heeejK-  ]r^-  (ju*  ]r_-  (jw*  ]r`-  (jy*  ]ra-  (hh	e]rb-  (hh	e]rc-  (hjN  e]rd-  (j~*  ]re-  (hhe]rf-  (hhe]rg-  (hjN  e]rh-  (j�*  ]ri-  (hh	e]rj-  (hh	eeee]rk-  (hh&ee]rl-  (h]rm-  (hh e]rn-  (hhe]ro-  (hhe]rp-  (h%heee]rq-  (ju*  ]rr-  (jw*  ]rs-  (jy*  ]rt-  (hh	e]ru-  (hh	e]rv-  (hjN  e]rw-  (j~*  ]rx-  (hhe]ry-  (hhe]rz-  (hjN  e]r{-  (j�*  ]r|-  (hh	e]r}-  (hh	eeee]r~-  (hh&ee]r-  (h]r�-  (hh e]r�-  (hhe]r�-  (hhe]r�-  (h%heee]r�-  (ju*  ]r�-  (jw*  ]r�-  (jy*  ]r�-  (hh	e]r�-  (hh	e]r�-  (hjN  e]r�-  (j~*  ]r�-  (hhe]r�-  (hhe]r�-  (hjN  e]r�-  (X	   Next-Mover�-  ]r�-  (hh	e]r�-  (hh	eeee]r�-  (hh&ee]r�-  (h]r�-  (hh e]r�-  (hhe]r�-  (hhe]r�-  (h%heee]r�-  (ju*  ]r�-  (jw*  ]r�-  (jy*  ]r�-  (hh	e]r�-  (hh	e]r�-  (hjN  e]r�-  (j~*  ]r�-  (hhe]r�-  (hhe]r�-  (hjN  e]r�-  (j�-  ]r�-  (hh	e]r�-  (hh	eeee]r�-  (hh&ee]r�-  (h]r�-  (hh e]r�-  (hhe]r�-  (hhe]r�-  (h%heeej�-  j�-  j�-  j�-  j�-  j�-  j�-  j�-  j�-  j�-  j�-  ]r�-  (ju*  ]r�-  (jw*  ]r�-  (jy*  ]r�-  (hh	e]r�-  (hh	e]r�-  (hjN  e]r�-  (j~*  ]r�-  (hhe]r�-  (hhe]r�-  (hjN  e]r�-  (j�-  ]r�-  (hh	e]r�-  (hh	eeee]r�-  (hh&ee]r�-  (h]r�-  (hh e]r�-  (hhe]r�-  (hhe]r�-  (h%heeej�-  ]r�-  (ju*  ]r�-  (jw*  ]r�-  (jy*  ]r�-  (hh	e]r�-  (hh	e]r�-  (hjN  e]r�-  (j~*  ]r�-  (hhe]r�-  (hhe]r�-  (hjN  e]r�-  (j�-  ]r�-  (hh	e]r�-  (hh	eeee]r�-  (hh&ee]r�-  (h]r�-  (hh e]r�-  (hhe]r�-  (hhe]r�-  (h%heeej�-  ]r�-  (ju*  ]r�-  (jw*  ]r�-  (jy*  ]r�-  (hh	e]r�-  (hh	e]r�-  (hjN  e]r�-  (j~*  ]r�-  (hhe]r�-  (hhe]r�-  (hjN  e]r�-  (j�-  ]r�-  (hh	e]r�-  (hh	eeee]r�-  (hh&ee]r�-  (h]r�-  (hh e]r�-  (hhe]r�-  (hhe]r�-  (h%heeej�-  j�-  j�-  ]r�-  (ju*  ]r�-  (jw*  ]r�-  (jy*  ]r�-  (hh	e]r�-  (hh	e]r�-  (hjN  e]r�-  (j~*  ]r�-  (hhe]r�-  (hhe]r�-  (hjN  e]r�-  (j�-  ]r�-  (hh	e]r�-  (hh	eeee]r�-  (hh&ee]r�-  (h]r�-  (hh e]r�-  (hhe]r�-  (hhe]r�-  (h%heeej�-  ]r�-  (ju*  ]r�-  (jw*  ]r�-  (jy*  ]r�-  (hh	e]r�-  (hh	e]r�-  (hjN  e]r�-  (j~*  ]r�-  (hhe]r�-  (hhe]r .  (hjN  e]r.  (j�-  ]r.  (hh	e]r.  (hh	eeee]r.  (hh&ee]r.  (h]r.  (hh e]r.  (hhe]r.  (hhe]r	.  (h%heee]r
.  (ju*  ]r.  (jw*  ]r.  (jy*  ]r.  (hh	e]r.  (hh	e]r.  (hjN  e]r.  (j~*  ]r.  (hhe]r.  (hhe]r.  (hjN  e]r.  (j�-  ]r.  (hh	e]r.  (hh	eeee]r.  (hh&ee]r.  (h]r.  (hh e]r.  (hhe]r.  (hhe]r.  (h%heeej
.  j
.  j
.  j
.  ]r.  (ju*  ]r.  (jw*  ]r.  (jy*  ]r .  (hh	e]r!.  (hh	e]r".  (hjN  e]r#.  (j~*  ]r$.  (hhe]r%.  (hhe]r&.  (hjN  e]r'.  (j�-  ]r(.  (hh	e]r).  (hh	eeee]r*.  (hh&ee]r+.  (h]r,.  (hh e]r-.  (hhe]r..  (hhe]r/.  (h%heeej.  j.  j.  ]r0.  (ju*  ]r1.  (jw*  ]r2.  (jy*  ]r3.  (hh	e]r4.  (hh	e]r5.  (hjN  e]r6.  (j~*  ]r7.  (hhe]r8.  (hhe]r9.  (hjN  e]r:.  (j�-  ]r;.  (hh	e]r<.  (hh	eeee]r=.  (hh&ee]r>.  (h]r?.  (hh e]r@.  (hhe]rA.  (hhe]rB.  (h%heeej0.  j0.  j0.  j0.  j0.  j0.  ]rC.  (ju*  ]rD.  (jw*  ]rE.  (jy*  ]rF.  (hh	e]rG.  (hh	e]rH.  (hjN  e]rI.  (j~*  ]rJ.  (hhe]rK.  (hhe]rL.  (hjN  e]rM.  (j�-  ]rN.  (hh	e]rO.  (hh	eeee]rP.  (hh&ee]rQ.  (h]rR.  (hh e]rS.  (hhe]rT.  (hhe]rU.  (h%heeejC.  jC.  jC.  ]rV.  (ju*  ]rW.  (jw*  ]rX.  (jy*  ]rY.  (hh	e]rZ.  (hh	e]r[.  (hjN  e]r\.  (j~*  ]r].  (hhe]r^.  (hhe]r_.  (hjN  e]r`.  (j�-  ]ra.  (hh	e]rb.  (hh	eeee]rc.  (hh&ee]rd.  (h]re.  (hh e]rf.  (hhe]rg.  (hhe]rh.  (h%heee]ri.  (ju*  ]rj.  (jw*  ]rk.  (jy*  ]rl.  (hh	e]rm.  (hh	e]rn.  (hjN  e]ro.  (j~*  ]rp.  (hhe]rq.  (hhe]rr.  (hjN  e]rs.  (j�-  ]rt.  (hh	e]ru.  (hh	eeee]rv.  (hh&ee]rw.  (h]rx.  (hh e]ry.  (hhe]rz.  (hhe]r{.  (h%heeeji.  ji.  ]r|.  (ju*  ]r}.  (jw*  ]r~.  (jy*  ]r.  (hh	e]r�.  (hh	e]r�.  (hjN  e]r�.  (j~*  ]r�.  (hhe]r�.  (hhe]r�.  (hjN  e]r�.  (j�-  ]r�.  (hh	e]r�.  (hh	eeee]r�.  (hh&ee]r�.  (h]r�.  (hh e]r�.  (hhe]r�.  (hhe]r�.  (h%heeej|.  ]r�.  (ju*  ]r�.  (jw*  ]r�.  (jy*  ]r�.  (hh	e]r�.  (hh	e]r�.  (hjN  e]r�.  (j~*  ]r�.  (hhe]r�.  (hhe]r�.  (hjN  e]r�.  (j�-  ]r�.  (hh	e]r�.  (hh	eeee]r�.  (hh&ee]r�.  (h]r�.  (hh e]r�.  (hhe]r�.  (hhe]r�.  (h%heeej�.  j�.  j�.  j�.  j�.  j�.  j�.  j�.  ]r�.  (ju*  ]r�.  (jw*  ]r�.  (jy*  ]r�.  (hh	e]r�.  (hh	e]r�.  (hjN  e]r�.  (j~*  ]r�.  (hhe]r�.  (hhe]r�.  (hjN  e]r�.  (j�-  ]r�.  (hh	e]r�.  (hh	eeee]r�.  (hh&ee]r�.  (h]r�.  (hh e]r�.  (hhe]r�.  (hhe]r�.  (h%heeej�.  ]r�.  (ju*  ]r�.  (jw*  ]r�.  (jy*  ]r�.  (hh	e]r�.  (hh	e]r�.  (hjN  e]r�.  (j~*  ]r�.  (hhe]r�.  (hhe]r�.  (hjN  e]r�.  (j�-  ]r�.  (hh	e]r�.  (hh	eeee]r�.  (hh&ee]r�.  (h]r�.  (hh e]r�.  (hhe]r�.  (hhe]r�.  (h%heee]r�.  (ju*  ]r�.  (jw*  ]r�.  (jy*  ]r�.  (hh	e]r�.  (hh	e]r�.  (hjN  e]r�.  (j~*  ]r�.  (hhe]r�.  (hhe]r�.  (hjN  e]r�.  (j�-  ]r�.  (hh	e]r�.  (hh	eeee]r�.  (hh&ee]r�.  (h]r�.  (hh e]r�.  (hhe]r�.  (hhe]r�.  (h%heeej�.  j�.  ]r�.  (ju*  ]r�.  (jw*  ]r�.  (jy*  ]r�.  (hh	e]r�.  (hh	e]r�.  (hjN  e]r�.  (j~*  ]r�.  (hhe]r�.  (hhe]r�.  (hjN  e]r�.  (j�-  ]r�.  (hh	e]r�.  (hh	eeee]r�.  (hh&ee]r�.  (h]r�.  (hh e]r�.  (hhe]r�.  (hhe]r�.  (h%heeej�.  j�.  ]r�.  (ju*  ]r�.  (jw*  ]r�.  (jy*  ]r�.  (hh	e]r�.  (hh	e]r�.  (hjN  e]r�.  (j~*  ]r�.  (hhe]r�.  (hhe]r�.  (hjN  e]r�.  (j�-  ]r�.  (hh	e]r�.  (hh	eeee]r�.  (hh&ee]r�.  (h]r�.  (hh e]r�.  (hhe]r�.  (hhe]r /  (h%heeej�.  ]r/  (ju*  ]r/  (jw*  ]r/  (jy*  ]r/  (hh	e]r/  (hh	e]r/  (hjN  e]r/  (j~*  ]r/  (hhe]r	/  (hhe]r
/  (hjN  e]r/  (j�-  ]r/  (hh	e]r/  (hh	eeee]r/  (hh&ee]r/  (h]r/  (hh e]r/  (hhe]r/  (hhe]r/  (h%heeej/  j/  j/  j/  ]r/  (ju*  ]r/  (jw*  ]r/  (jy*  ]r/  (hh	e]r/  (hh	e]r/  (hjN  e]r/  (j~*  ]r/  (hhe]r/  (hhe]r/  (hjN  e]r/  (j�-  ]r/  (hh	e]r /  (hh	eeee]r!/  (hh&ee]r"/  (h]r#/  (hh e]r$/  (hhe]r%/  (hhe]r&/  (h%heeej/  j/  j/  j/  j/  j/  j/  j/  j/  ]r'/  (ju*  ]r(/  (jw*  ]r)/  (jy*  ]r*/  (hh	e]r+/  (hh	e]r,/  (hjN  e]r-/  (j~*  ]r./  (hhe]r//  (hhe]r0/  (hjN  e]r1/  (j�-  ]r2/  (hh	e]r3/  (hh	eeee]r4/  (hh&ee]r5/  (h]r6/  (hh e]r7/  (hhe]r8/  (hhe]r9/  (h%heeej'/  j'/  j'/  j'/  j'/  j'/  j'/  j'/  ]r:/  (ju*  ]r;/  (jw*  ]r</  (jy*  ]r=/  (hh	e]r>/  (hh	e]r?/  (hjN  e]r@/  (j~*  ]rA/  (hhe]rB/  (hhe]rC/  (hjN  e]rD/  (j�-  ]rE/  (hh	e]rF/  (hh	eeee]rG/  (hh&ee]rH/  (h]rI/  (hh e]rJ/  (hhe]rK/  (hhe]rL/  (h%heee]rM/  (ju*  ]rN/  (jw*  ]rO/  (jy*  ]rP/  (hh	e]rQ/  (hh	e]rR/  (hjN  e]rS/  (j~*  ]rT/  (hhe]rU/  (hhe]rV/  (hjN  e]rW/  (j�-  ]rX/  (hh	e]rY/  (hh	eeee]rZ/  (hh&ee]r[/  (h]r\/  (hh e]r]/  (hhe]r^/  (hhe]r_/  (h%heeejM/  jM/  jM/  jM/  jM/  jM/  jM/  jM/  ]r`/  (ju*  ]ra/  (jw*  ]rb/  (jy*  ]rc/  (hh	e]rd/  (hh	e]re/  (hjN  e]rf/  (j~*  ]rg/  (hhe]rh/  (hhe]ri/  (hjN  e]rj/  (j�-  ]rk/  (hh	e]rl/  (hh	eeee]rm/  (hh&ee]rn/  (h]ro/  (hh e]rp/  (hhe]rq/  (hhe]rr/  (h%heeej`/  j`/  j`/  j`/  j`/  j`/  j`/  j`/  ]rs/  (ju*  ]rt/  (jw*  ]ru/  (jy*  ]rv/  (hh	e]rw/  (hh	e]rx/  (hjN  e]ry/  (j~*  ]rz/  (hhe]r{/  (hhe]r|/  (hjN  e]r}/  (j�-  ]r~/  (hh	e]r/  (hh	eeee]r�/  (hh&ee]r�/  (h]r�/  (hh e]r�/  (hhe]r�/  (hhe]r�/  (h%heeejs/  js/  js/  js/  js/  js/  ]r�/  (ju*  ]r�/  (jw*  ]r�/  (jy*  ]r�/  (hh	e]r�/  (hh	e]r�/  (hjN  e]r�/  (j~*  ]r�/  (hhe]r�/  (hhe]r�/  (hjN  e]r�/  (j�-  ]r�/  (hh	e]r�/  (hh	eeee]r�/  (hh&ee]r�/  (h]r�/  (hh e]r�/  (hhe]r�/  (hhe]r�/  (h%heee]r�/  (ju*  ]r�/  (jw*  ]r�/  (jy*  ]r�/  (hh	e]r�/  (hh	e]r�/  (hjN  e]r�/  (j~*  ]r�/  (hhe]r�/  (hhe]r�/  (hjN  e]r�/  (j�-  ]r�/  (hh	e]r�/  (hh	eeee]r�/  (hh&ee]r�/  (h]r�/  (hh e]r�/  (hhe]r�/  (hhe]r�/  (h%heee]r�/  (ju*  ]r�/  (jw*  ]r�/  (jy*  ]r�/  (hh	e]r�/  (hh	e]r�/  (hjN  e]r�/  (j~*  ]r�/  (hhe]r�/  (hhe]r�/  (hjN  e]r�/  (j�-  ]r�/  (hh	e]r�/  (hh	eeee]r�/  (hh&ee]r�/  (h]r�/  (hh e]r�/  (hhe]r�/  (hhe]r�/  (h%heeej�/  j�/  j�/  j�/  ]r�/  (ju*  ]r�/  (jw*  ]r�/  (jy*  ]r�/  (hh	e]r�/  (hh	e]r�/  (hjN  e]r�/  (j~*  ]r�/  (hhe]r�/  (hhe]r�/  (hjN  e]r�/  (j�-  ]r�/  (hh	e]r�/  (hh	eeee]r�/  (hh&ee]r�/  (h]r�/  (hh e]r�/  (hhe]r�/  (hhe]r�/  (h%heeej�/  ]r�/  (ju*  ]r�/  (jw*  ]r�/  (jy*  ]r�/  (hh	e]r�/  (hh	e]r�/  (hjN  e]r�/  (j~*  ]r�/  (hhe]r�/  (hhe]r�/  (hjN  e]r�/  (j�-  ]r�/  (hh	e]r�/  (hh	eeee]r�/  (hh&ee]r�/  (h]r�/  (hh e]r�/  (hhe]r�/  (hhe]r�/  (h%heeej�/  j�/  ]r�/  (ju*  ]r�/  (jw*  ]r�/  (jy*  ]r�/  (hh	e]r�/  (hh	e]r�/  (hjN  e]r�/  (j~*  ]r�/  (hhe]r�/  (hhe]r�/  (hjN  e]r�/  (j�-  ]r�/  (hh	e]r�/  (hh	eeee]r�/  (hh&ee]r�/  (h]r�/  (hh e]r�/  (hhe]r�/  (hhe]r�/  (h%heeej�/  j�/  j�/  j�/  j�/  j�/  j�/  ]r�/  (ju*  ]r�/  (jw*  ]r�/  (jy*  ]r�/  (hh	e]r�/  (hh	e]r�/  (hjN  e]r�/  (j~*  ]r�/  (hhe]r 0  (hhe]r0  (hjN  e]r0  (j�-  ]r0  (hh	e]r0  (hh	eeee]r0  (hh&ee]r0  (h]r0  (hh e]r0  (hhe]r	0  (hhe]r
0  (h%heeej�/  j�/  ]r0  (ju*  ]r0  (jw*  ]r0  (jy*  ]r0  (hh	e]r0  (hh	e]r0  (hjN  e]r0  (j~*  ]r0  (hhe]r0  (hhe]r0  (hjN  e]r0  (j�-  ]r0  (hh	e]r0  (hh	eeee]r0  (hh&ee]r0  (h]r0  (hh e]r0  (hhe]r0  (hhe]r0  (h%heeej0  j0  j0  ]r0  (ju*  ]r0  (jw*  ]r 0  (jy*  ]r!0  (hh	e]r"0  (hh	e]r#0  (hjN  e]r$0  (j~*  ]r%0  (hhe]r&0  (hhe]r'0  (hjN  e]r(0  (j�-  ]r)0  (hh	e]r*0  (hh	eeee]r+0  (hh&ee]r,0  (h]r-0  (hh e]r.0  (hhe]r/0  (hhe]r00  (h%heeej0  j0  ]r10  (ju*  ]r20  (jw*  ]r30  (jy*  ]r40  (hh	e]r50  (hh	e]r60  (hjN  e]r70  (j~*  ]r80  (hhe]r90  (hhe]r:0  (hjN  e]r;0  (j�-  ]r<0  (hh	e]r=0  (hh	eeee]r>0  (hh&ee]r?0  (h]r@0  (hh e]rA0  (hhe]rB0  (hhe]rC0  (h%heeej10  j10  ]rD0  (ju*  ]rE0  (jw*  ]rF0  (jy*  ]rG0  (hh	e]rH0  (hh	e]rI0  (hjN  e]rJ0  (j~*  ]rK0  (hhe]rL0  (hhe]rM0  (hjN  e]rN0  (j�-  ]rO0  (hh	e]rP0  (hh	eeee]rQ0  (hh&ee]rR0  (h]rS0  (hh e]rT0  (hhe]rU0  (hhe]rV0  (h%heeejD0  jD0  ]rW0  (ju*  ]rX0  (jw*  ]rY0  (jy*  ]rZ0  (hh	e]r[0  (hh	e]r\0  (hjN  e]r]0  (j~*  ]r^0  (hhe]r_0  (hhe]r`0  (hjN  e]ra0  (j�-  ]rb0  (hh	e]rc0  (hh	eeee]rd0  (hh&ee]re0  (h]rf0  (hh e]rg0  (hhe]rh0  (hhe]ri0  (h%heeejW0  ]rj0  (ju*  ]rk0  (jw*  ]rl0  (jy*  ]rm0  (hh	e]rn0  (hh	e]ro0  (hjN  e]rp0  (j~*  ]rq0  (hhe]rr0  (hhe]rs0  (hjN  e]rt0  (j�-  ]ru0  (hh	e]rv0  (hh	eeee]rw0  (hh&ee]rx0  (h]ry0  (hh e]rz0  (hhe]r{0  (hhe]r|0  (h%heeejj0  jj0  jj0  ]r}0  (ju*  ]r~0  (jw*  ]r0  (jy*  ]r�0  (hh	e]r�0  (hh	e]r�0  (hjN  e]r�0  (j~*  ]r�0  (hhe]r�0  (hhe]r�0  (hjN  e]r�0  (j�-  ]r�0  (hh	e]r�0  (hh	eeee]r�0  (hh&ee]r�0  (h]r�0  (hh e]r�0  (hhe]r�0  (hhe]r�0  (h%heeej}0  j}0  j}0  ]r�0  (ju*  ]r�0  (jw*  ]r�0  (jy*  ]r�0  (hh	e]r�0  (hh	e]r�0  (hjN  e]r�0  (j~*  ]r�0  (hhe]r�0  (hhe]r�0  (hjN  e]r�0  (j�-  ]r�0  (hh	e]r�0  (hh	eeee]r�0  (hh&ee]r�0  (h]r�0  (hh e]r�0  (hhe]r�0  (hhe]r�0  (h%heeej�0  j�0  j�0  ]r�0  (ju*  ]r�0  (jw*  ]r�0  (jy*  ]r�0  (hh	e]r�0  (hh	e]r�0  (hjN  e]r�0  (j~*  ]r�0  (hhe]r�0  (hhe]r�0  (hjN  e]r�0  (j�-  ]r�0  (hh	e]r�0  (hh	eeee]r�0  (hh&ee]r�0  (h]r�0  (hh e]r�0  (hhe]r�0  (hhe]r�0  (h%heeej�0  ]r�0  (ju*  ]r�0  (jw*  ]r�0  (jy*  ]r�0  (hh	e]r�0  (hh	e]r�0  (hjN  e]r�0  (j~*  ]r�0  (hhe]r�0  (hhe]r�0  (hjN  e]r�0  (j�-  ]r�0  (hh	e]r�0  (hh	eeee]r�0  (hh&ee]r�0  (h]r�0  (hh e]r�0  (hhe]r�0  (hhe]r�0  (h%heeej�0  j�0  j�0  j�0  ]r�0  (ju*  ]r�0  (jw*  ]r�0  (jy*  ]r�0  (hh	e]r�0  (hh	e]r�0  (hjN  e]r�0  (j~*  ]r�0  (hhe]r�0  (hhe]r�0  (hjN  e]r�0  (j�-  ]r�0  (hh	e]r�0  (hh	eeee]r�0  (hh&ee]r�0  (h]r�0  (hh e]r�0  (hhe]r�0  (hhe]r�0  (h%heeej�0  ]r�0  (ju*  ]r�0  (jw*  ]r�0  (jy*  ]r�0  (hh	e]r�0  (hh	e]r�0  (hjN  e]r�0  (j~*  ]r�0  (hhe]r�0  (hhe]r�0  (hjN  e]r�0  (j�-  ]r�0  (hh	e]r�0  (hh	eeee]r�0  (hh&ee]r�0  (h]r�0  (hh e]r�0  (hhe]r�0  (hhe]r�0  (h%heeej�0  ]r�0  (ju*  ]r�0  (jw*  ]r�0  (jy*  ]r�0  (hh	e]r�0  (hh	e]r�0  (hjN  e]r�0  (j~*  ]r�0  (hhe]r�0  (hhe]r�0  (hjN  e]r�0  (j�-  ]r�0  (hh	e]r�0  (hh	eeee]r�0  (hh&ee]r�0  (h]r�0  (hh e]r�0  (hhe]r 1  (hhe]r1  (h%heeej�0  j�0  j�0  ]r1  (ju*  ]r1  (jw*  ]r1  (jy*  ]r1  (hh	e]r1  (hh	e]r1  (hjN  e]r1  (j~*  ]r	1  (hh	e]r
1  (hhe]r1  (hjN  e]r1  (j�-  ]r1  (hh	e]r1  (hh	eeee]r1  (hh&ee]r1  (h]r1  (hh e]r1  (hhe]r1  (hhe]r1  (h%heeej1  ]r1  (ju*  ]r1  (jw*  ]r1  (jy*  ]r1  (hh	e]r1  (hh	e]r1  (hjN  e]r1  (j~*  ]r1  (hh	e]r1  (hhe]r1  (hjN  e]r1  (j�-  ]r 1  (hh	e]r!1  (hh	eeee]r"1  (hh&ee]r#1  (h]r$1  (hh e]r%1  (hhe]r&1  (hhe]r'1  (h%heeej1  j1  j1  ]r(1  (ju*  ]r)1  (jw*  ]r*1  (jy*  ]r+1  (hh	e]r,1  (hh	e]r-1  (hjN  e]r.1  (j~*  ]r/1  (hh	e]r01  (hhe]r11  (hjN  e]r21  (j�-  ]r31  (hh	e]r41  (hh	eeee]r51  (hh&ee]r61  (h]r71  (hh e]r81  (hhe]r91  (hhe]r:1  (h%heeej(1  j(1  j(1  j(1  ]r;1  (ju*  ]r<1  (jw*  ]r=1  (jy*  ]r>1  (hh	e]r?1  (hh	e]r@1  (hjN  e]rA1  (j~*  ]rB1  (hh	e]rC1  (hhe]rD1  (hjN  e]rE1  (j�-  ]rF1  (hh	e]rG1  (hh	eeee]rH1  (hh&ee]rI1  (h]rJ1  (hh e]rK1  (hhe]rL1  (hhe]rM1  (h%heeej;1  j;1  ]rN1  (ju*  ]rO1  (jw*  ]rP1  (jy*  ]rQ1  (hh	e]rR1  (hh	e]rS1  (hjN  e]rT1  (j~*  ]rU1  (hh	e]rV1  (hhe]rW1  (hjN  e]rX1  (j�-  ]rY1  (hh	e]rZ1  (hh	eeee]r[1  (hh&ee]r\1  (h]r]1  (hh e]r^1  (hhe]r_1  (hhe]r`1  (h%heee]ra1  (ju*  ]rb1  (jw*  ]rc1  (jy*  ]rd1  (hh	e]re1  (hh	e]rf1  (hjN  e]rg1  (j~*  ]rh1  (hh	e]ri1  (hhe]rj1  (hjN  e]rk1  (j�-  ]rl1  (hh	e]rm1  (hh	eeee]rn1  (hh&ee]ro1  (h]rp1  (hh e]rq1  (hhe]rr1  (hhe]rs1  (h%heeeja1  ja1  ja1  ja1  ]rt1  (ju*  ]ru1  (jw*  ]rv1  (jy*  ]rw1  (hh	e]rx1  (hh	e]ry1  (hjN  e]rz1  (j~*  ]r{1  (hh	e]r|1  (hhe]r}1  (hjN  e]r~1  (j�-  ]r1  (hh	e]r�1  (hh	eeee]r�1  (hh&ee]r�1  (h]r�1  (hh e]r�1  (hhe]r�1  (hhe]r�1  (h%heeejt1  ]r�1  (ju*  ]r�1  (jw*  ]r�1  (jy*  ]r�1  (hh	e]r�1  (hh	e]r�1  (hjN  e]r�1  (j~*  ]r�1  (hhe]r�1  (hhe]r�1  (hjN  e]r�1  (j�-  ]r�1  (hh	e]r�1  (hh	eeee]r�1  (hh&ee]r�1  (h]r�1  (hh e]r�1  (hhe]r�1  (hhe]r�1  (h%heeej�1  ]r�1  (ju*  ]r�1  (jw*  ]r�1  (jy*  ]r�1  (hh	e]r�1  (hh	e]r�1  (hjN  e]r�1  (j~*  ]r�1  (hhe]r�1  (hhe]r�1  (hjN  e]r�1  (j�-  ]r�1  (hh	e]r�1  (hh	eeee]r�1  (hh&ee]r�1  (h]r�1  (hh e]r�1  (hhe]r�1  (hhe]r�1  (h%heeej�1  j�1  j�1  ]r�1  (ju*  ]r�1  (jw*  ]r�1  (jy*  ]r�1  (hh	e]r�1  (hh	e]r�1  (hjN  e]r�1  (j~*  ]r�1  (hhe]r�1  (hhe]r�1  (hjN  e]r�1  (j�-  ]r�1  (hh	e]r�1  (hh	eeee]r�1  (hh&ee]r�1  (h]r�1  (hh e]r�1  (hhe]r�1  (hhe]r�1  (h%heeej�1  j�1  j�1  j�1  j�1  j�1  j�1  j�1  ]r�1  (ju*  ]r�1  (jw*  ]r�1  (jy*  ]r�1  (hh	e]r�1  (hh	e]r�1  (hjN  e]r�1  (j~*  ]r�1  (hhe]r�1  (hhe]r�1  (hjN  e]r�1  (j�-  ]r�1  (hh	e]r�1  (hh	eeee]r�1  (hh&ee]r�1  (h]r�1  (hh e]r�1  (hhe]r�1  (hhe]r�1  (h%heee]r�1  (ju*  ]r�1  (jw*  ]r�1  (jy*  ]r�1  (hh	e]r�1  (hh	e]r�1  (hjN  e]r�1  (j~*  ]r�1  (hhe]r�1  (hhe]r�1  (hjN  e]r�1  (j�-  ]r�1  (hh	e]r�1  (hh	eeee]r�1  (hh&ee]r�1  (h]r�1  (hh e]r�1  (hhe]r�1  (hhe]r�1  (h%heee]r�1  (ju*  ]r�1  (jw*  ]r�1  (jy*  ]r�1  (hh	e]r�1  (hh	e]r�1  (hjN  e]r�1  (j~*  ]r�1  (hhe]r�1  (hhe]r�1  (hjN  e]r�1  (j�-  ]r�1  (hh	e]r�1  (hh	eeee]r�1  (hh&ee]r�1  (h]r�1  (hh e]r�1  (hhe]r�1  (hhe]r�1  (h%heeej�1  j�1  ]r�1  (ju*  ]r�1  (jw*  ]r�1  (jy*  ]r�1  (hh	e]r�1  (hh	e]r�1  (hjN  e]r�1  (j~*  ]r 2  (hhe]r2  (hhe]r2  (hjN  e]r2  (j�-  ]r2  (hh	e]r2  (hh	eeee]r2  (hh&ee]r2  (h]r2  (hh e]r	2  (hhe]r
2  (hhe]r2  (h%heeej�1  ]r2  (ju*  ]r2  (jw*  ]r2  (jy*  ]r2  (hh	e]r2  (hh	e]r2  (hjN  e]r2  (j~*  ]r2  (hhe]r2  (hhe]r2  (hjN  e]r2  (j�-  ]r2  (hh	e]r2  (hh	eeee]r2  (hh&ee]r2  (h]r2  (hh e]r2  (hhe]r2  (hhe]r2  (h%heeej2  ]r2  (ju*  ]r 2  (jw*  ]r!2  (jy*  ]r"2  (hh	e]r#2  (hh	e]r$2  (hjN  e]r%2  (j~*  ]r&2  (hhe]r'2  (hhe]r(2  (hjN  e]r)2  (j�-  ]r*2  (hh	e]r+2  (hh	eeee]r,2  (hh&ee]r-2  (h]r.2  (hh e]r/2  (hhe]r02  (hhe]r12  (h%heeej2  j2  ]r22  (ju*  ]r32  (jw*  ]r42  (jy*  ]r52  (hh	e]r62  (hh	e]r72  (hjN  e]r82  (j~*  ]r92  (hhe]r:2  (hhe]r;2  (hjN  e]r<2  (j�-  ]r=2  (hh	e]r>2  (hh	eeee]r?2  (hh&ee]r@2  (h]rA2  (hh e]rB2  (hhe]rC2  (hhe]rD2  (h%heeej22  j22  j22  j22  j22  j22  ]rE2  (ju*  ]rF2  (jw*  ]rG2  (jy*  ]rH2  (hh	e]rI2  (hh	e]rJ2  (hjN  e]rK2  (j~*  ]rL2  (hhe]rM2  (hhe]rN2  (hjN  e]rO2  (j�-  ]rP2  (hh	e]rQ2  (hh	eeee]rR2  (hh&ee]rS2  (h]rT2  (hh e]rU2  (hhe]rV2  (hh	e]rW2  (h%heeejE2  jE2  ]rX2  (ju*  ]rY2  (jw*  ]rZ2  (jy*  ]r[2  (hh	e]r\2  (hh	e]r]2  (hjN  e]r^2  (j~*  ]r_2  (hhe]r`2  (hhe]ra2  (hjN  e]rb2  (j�-  ]rc2  (hh	e]rd2  (hh	eeee]re2  (hh&ee]rf2  (h]rg2  (hh e]rh2  (hhe]ri2  (hh	e]rj2  (h%heee]rk2  (ju*  ]rl2  (jw*  ]rm2  (jy*  ]rn2  (hh	e]ro2  (hh	e]rp2  (hjN  e]rq2  (j~*  ]rr2  (hhe]rs2  (hhe]rt2  (hjN  e]ru2  (j�-  ]rv2  (hh	e]rw2  (hh	eeee]rx2  (hh&ee]ry2  (h]rz2  (hh e]r{2  (hhe]r|2  (hhe]r}2  (h%heeejk2  jk2  jk2  jk2  jk2  ]r~2  (ju*  ]r2  (jw*  ]r�2  (jy*  ]r�2  (hh	e]r�2  (hh	e]r�2  (hjN  e]r�2  (j~*  ]r�2  (hhe]r�2  (hhe]r�2  (hjN  e]r�2  (j�-  ]r�2  (hh	e]r�2  (hh	eeee]r�2  (hh&ee]r�2  (h]r�2  (hh e]r�2  (hhe]r�2  (hhe]r�2  (h%heee]r�2  (ju*  ]r�2  (jw*  ]r�2  (jy*  ]r�2  (hh	e]r�2  (hh	e]r�2  (hjN  e]r�2  (j~*  ]r�2  (hhe]r�2  (hhe]r�2  (hjN  e]r�2  (j�-  ]r�2  (hh	e]r�2  (hh	eeee]r�2  (hh&ee]r�2  (h]r�2  (hh e]r�2  (hhe]r�2  (hhe]r�2  (h%heee]r�2  (ju*  ]r�2  (jw*  ]r�2  (jy*  ]r�2  (hh	e]r�2  (hh	e]r�2  (hjN  e]r�2  (j~*  ]r�2  (hhe]r�2  (hhe]r�2  (hjN  e]r�2  (j�-  ]r�2  (hh	e]r�2  (hh	eeee]r�2  (hh&ee]r�2  (h]r�2  (hh e]r�2  (hhe]r�2  (hhe]r�2  (h%heee]r�2  (ju*  ]r�2  (jw*  ]r�2  (jy*  ]r�2  (hh	e]r�2  (hh	e]r�2  (hjN  e]r�2  (j~*  ]r�2  (hhe]r�2  (hhe]r�2  (hjN  e]r�2  (j�-  ]r�2  (hh	e]r�2  (hh	eeee]r�2  (hh&ee]r�2  (h]r�2  (hh e]r�2  (hhe]r�2  (hhe]r�2  (h%heeej�2  j�2  j�2  j�2  j�2  ]r�2  (ju*  ]r�2  (jw*  ]r�2  (jy*  ]r�2  (hh	e]r�2  (hh	e]r�2  (hjN  e]r�2  (j~*  ]r�2  (hhe]r�2  (hhe]r�2  (hjN  e]r�2  (j�-  ]r�2  (hh	e]r�2  (hh	eeee]r�2  (hh&ee]r�2  (h]r�2  (hh e]r�2  (hhe]r�2  (hhe]r�2  (h%heeej�2  j�2  j�2  j�2  j�2  j�2  j�2  ]r�2  (ju*  ]r�2  (jw*  ]r�2  (jy*  ]r�2  (hh	e]r�2  (hh	e]r�2  (hjN  e]r�2  (j~*  ]r�2  (hhe]r�2  (hhe]r�2  (hjN  e]r�2  (j�-  ]r�2  (hh	e]r�2  (hh	eeee]r�2  (hh&ee]r�2  (h]r�2  (hh e]r�2  (hhe]r�2  (hhe]r�2  (h%heeej�2  j�2  j�2  j�2  ]r�2  (ju*  ]r�2  (jw*  ]r�2  (jy*  ]r�2  (hh	e]r�2  (hh	e]r�2  (hjN  e]r�2  (j~*  ]r�2  (hhe]r�2  (hhe]r�2  (hjN  e]r�2  (j�-  ]r�2  (hh	e]r�2  (hh	eeee]r�2  (hh&ee]r�2  (h]r�2  (hh e]r 3  (hhe]r3  (hhe]r3  (h%heeej�2  ]r3  (ju*  ]r3  (jw*  ]r3  (jy*  ]r3  (hh	e]r3  (hh	e]r3  (hjN  e]r	3  (j~*  ]r
3  (hhe]r3  (hhe]r3  (hjN  e]r3  (j�-  ]r3  (hh	e]r3  (hh	eeee]r3  (hh&ee]r3  (h]r3  (hh e]r3  (hhe]r3  (hhe]r3  (h%heeej3  j3  j3  j3  j3  j3  j3  j3  j3  j3  ]r3  (ju*  ]r3  (jw*  ]r3  (jy*  ]r3  (hh	e]r3  (hh	e]r3  (hjN  e]r3  (j~*  ]r3  (hhe]r3  (hhe]r3  (hjN  e]r 3  (j�-  ]r!3  (hh	e]r"3  (hh	eeee]r#3  (hh&ee]r$3  (h]r%3  (hh e]r&3  (hhe]r'3  (hhe]r(3  (h%heeej3  j3  j3  j3  j3  j3  j3  j3  j3  j3  ]r)3  (ju*  ]r*3  (jw*  ]r+3  (jy*  ]r,3  (hh	e]r-3  (hh	e]r.3  (hjN  e]r/3  (j~*  ]r03  (hhe]r13  (hhe]r23  (hjN  e]r33  (j�-  ]r43  (hh	e]r53  (hh	eeee]r63  (hh&ee]r73  (h]r83  (hh e]r93  (hhe]r:3  (hhe]r;3  (h%heee]r<3  (ju*  ]r=3  (jw*  ]r>3  (jy*  ]r?3  (hh	e]r@3  (hh	e]rA3  (hjN  e]rB3  (j~*  ]rC3  (hhe]rD3  (hhe]rE3  (hjN  e]rF3  (j�-  ]rG3  (hh	e]rH3  (hh	eeee]rI3  (hh&ee]rJ3  (h]rK3  (hh e]rL3  (hhe]rM3  (hhe]rN3  (h%heeej<3  j<3  j<3  j<3  j<3  j<3  j<3  j<3  j<3  j<3  j<3  j<3  j<3  ]rO3  (ju*  ]rP3  (jw*  ]rQ3  (jy*  ]rR3  (hh	e]rS3  (hh	e]rT3  (hjN  e]rU3  (j~*  ]rV3  (hhe]rW3  (hhe]rX3  (hjN  e]rY3  (j�-  ]rZ3  (hh	e]r[3  (hh	eeee]r\3  (hh&ee]r]3  (h]r^3  (hh e]r_3  (hhe]r`3  (hhe]ra3  (h%heee]rb3  (ju*  ]rc3  (jw*  ]rd3  (jy*  ]re3  (hh	e]rf3  (hh	e]rg3  (hjN  e]rh3  (j~*  ]ri3  (hhe]rj3  (hhe]rk3  (hjN  e]rl3  (j�-  ]rm3  (hh	e]rn3  (hh	eeee]ro3  (hh&ee]rp3  (h]rq3  (hh e]rr3  (hhe]rs3  (hhe]rt3  (h%heee]ru3  (ju*  ]rv3  (jw*  ]rw3  (jy*  ]rx3  (hh	e]ry3  (hh	e]rz3  (hjN  e]r{3  (j~*  ]r|3  (hhe]r}3  (hhe]r~3  (hjN  e]r3  (j�-  ]r�3  (hh	e]r�3  (hh	eeee]r�3  (hh&ee]r�3  (h]r�3  (hh e]r�3  (hhe]r�3  (hhe]r�3  (h%heeeju3  ]r�3  (ju*  ]r�3  (jw*  ]r�3  (jy*  ]r�3  (hh	e]r�3  (hh	e]r�3  (hjN  e]r�3  (j~*  ]r�3  (hhe]r�3  (hhe]r�3  (hjN  e]r�3  (j�-  ]r�3  (hh	e]r�3  (hh	eeee]r�3  (hh&ee]r�3  (h]r�3  (hh e]r�3  (hhe]r�3  (hhe]r�3  (h%heee]r�3  (ju*  ]r�3  (jw*  ]r�3  (jy*  ]r�3  (hh	e]r�3  (hh	e]r�3  (hjN  e]r�3  (j~*  ]r�3  (hhe]r�3  (hhe]r�3  (hjN  e]r�3  (j�-  ]r�3  (hh	e]r�3  (hh	eeee]r�3  (hh&ee]r�3  (h]r�3  (hh e]r�3  (hhe]r�3  (hhe]r�3  (h%heee]r�3  (ju*  ]r�3  (jw*  ]r�3  (jy*  ]r�3  (hh	e]r�3  (hh	e]r�3  (hjN  e]r�3  (j~*  ]r�3  (hhe]r�3  (hhe]r�3  (hjN  e]r�3  (j�-  ]r�3  (hh	e]r�3  (hh	eeee]r�3  (hh&ee]r�3  (h]r�3  (hh e]r�3  (hhe]r�3  (hhe]r�3  (h%heeej�3  ]r�3  (ju*  ]r�3  (jw*  ]r�3  (jy*  ]r�3  (hh	e]r�3  (hh	e]r�3  (hjN  e]r�3  (j~*  ]r�3  (hh	e]r�3  (hhe]r�3  (hjN  e]r�3  (j�-  ]r�3  (hh	e]r�3  (hh	eeee]r�3  (hh&ee]r�3  (h]r�3  (hh e]r�3  (hhe]r�3  (hhe]r�3  (h%heee]r�3  (ju*  ]r�3  (jw*  ]r�3  (jy*  ]r�3  (hh	e]r�3  (hh	e]r�3  (hjN  e]r�3  (j~*  ]r�3  (hh	e]r�3  (hhe]r�3  (hjN  e]r�3  (j�-  ]r�3  (hh	e]r�3  (hh	eeee]r�3  (hh&ee]r�3  (h]r�3  (hh e]r�3  (hhe]r�3  (hhe]r�3  (h%heeej�3  j�3  j�3  j�3  ]r�3  (ju*  ]r�3  (jw*  ]r�3  (jy*  ]r�3  (hh	e]r�3  (hh	e]r�3  (hjN  e]r�3  (j~*  ]r�3  (hh	e]r�3  (hhe]r�3  (hjN  e]r�3  (j�-  ]r�3  (hh	e]r�3  (hh	eeee]r�3  (hh&ee]r�3  (h]r�3  (hh e]r�3  (hhe]r�3  (hhe]r�3  (h%heee]r�3  (ju*  ]r�3  (jw*  ]r�3  (jy*  ]r�3  (hh	e]r�3  (hh	e]r�3  (hjN  e]r 4  (j~*  ]r4  (hh	e]r4  (hhe]r4  (hjN  e]r4  (j�-  ]r4  (hh	e]r4  (hh	eeee]r4  (hh&ee]r4  (h]r	4  (hh e]r
4  (hhe]r4  (hhe]r4  (h%heeej�3  ]r4  (ju*  ]r4  (jw*  ]r4  (jy*  ]r4  (hh	e]r4  (hh	e]r4  (hjN  e]r4  (j~*  ]r4  (hh	e]r4  (hhe]r4  (hjN  e]r4  (j�-  ]r4  (hh	e]r4  (hh	eeee]r4  (hh&ee]r4  (h]r4  (hh e]r4  (hhe]r4  (hhe]r4  (h%heeej4  ]r 4  (ju*  ]r!4  (jw*  ]r"4  (jy*  ]r#4  (hh	e]r$4  (hh	e]r%4  (hjN  e]r&4  (j~*  ]r'4  (hh	e]r(4  (hhe]r)4  (hjN  e]r*4  (j�-  ]r+4  (hh	e]r,4  (hh	eeee]r-4  (hh&ee]r.4  (h]r/4  (hh e]r04  (hhe]r14  (hh	e]r24  (h%heeej 4  j 4  j 4  ]r34  (ju*  ]r44  (jw*  ]r54  (jy*  ]r64  (hh	e]r74  (hh	e]r84  (hjN  e]r94  (j~*  ]r:4  (hh	e]r;4  (hhe]r<4  (hjN  e]r=4  (j�-  ]r>4  (hh	e]r?4  (hh	eeee]r@4  (hh&ee]rA4  (h]rB4  (hh e]rC4  (hhe]rD4  (hh	e]rE4  (h%heeej34  j34  j34  j34  j34  j34  ]rF4  (ju*  ]rG4  (jw*  ]rH4  (jy*  ]rI4  (hh	e]rJ4  (hh	e]rK4  (hjN  e]rL4  (j~*  ]rM4  (hh	e]rN4  (hhe]rO4  (hjN  e]rP4  (j�-  ]rQ4  (hh	e]rR4  (hh	eeee]rS4  (hh&ee]rT4  (h]rU4  (hh e]rV4  (hhe]rW4  (hh	e]rX4  (h%heeejF4  jF4  ]rY4  (ju*  ]rZ4  (jw*  ]r[4  (jy*  ]r\4  (hh	e]r]4  (hh	e]r^4  (hjN  e]r_4  (j~*  ]r`4  (hh	e]ra4  (hhe]rb4  (hjN  e]rc4  (j�-  ]rd4  (hh	e]re4  (hh	eeee]rf4  (hh&ee]rg4  (h]rh4  (hh e]ri4  (hhe]rj4  (hh	e]rk4  (h%heeejY4  jY4  ]rl4  (ju*  ]rm4  (jw*  ]rn4  (jy*  ]ro4  (hh	e]rp4  (hh	e]rq4  (hjN  e]rr4  (j~*  ]rs4  (hh	e]rt4  (hhe]ru4  (hjN  e]rv4  (j�-  ]rw4  (hh	e]rx4  (hh	eeee]ry4  (hh&ee]rz4  (h]r{4  (hh e]r|4  (hhe]r}4  (hh	e]r~4  (h%heeejl4  ]r4  (ju*  ]r�4  (jw*  ]r�4  (jy*  ]r�4  (hh	e]r�4  (hh	e]r�4  (hjN  e]r�4  (j~*  ]r�4  (hh	e]r�4  (hhe]r�4  (hjN  e]r�4  (j�-  ]r�4  (hh	e]r�4  (hh	eeee]r�4  (hh&ee]r�4  (h]r�4  (hh e]r�4  (hhe]r�4  (hh	e]r�4  (h%heeej4  j4  j4  j4  ]r�4  (ju*  ]r�4  (jw*  ]r�4  (jy*  ]r�4  (hh	e]r�4  (hh	e]r�4  (hjN  e]r�4  (j~*  ]r�4  (hh	e]r�4  (hhe]r�4  (hjN  e]r�4  (j�-  ]r�4  (hh	e]r�4  (hh	eeee]r�4  (hh&ee]r�4  (h]r�4  (hh e]r�4  (hhe]r�4  (hh	e]r�4  (h%heee]r�4  (ju*  ]r�4  (jw*  ]r�4  (jy*  ]r�4  (hh	e]r�4  (hh	e]r�4  (hjN  e]r�4  (j~*  ]r�4  (hh	e]r�4  (hhe]r�4  (hjN  e]r�4  (j�-  ]r�4  (hh	e]r�4  (hh	eeee]r�4  (hh&ee]r�4  (h]r�4  (hh e]r�4  (hhe]r�4  (hh	e]r�4  (h%heeej�4  j�4  ]r�4  (ju*  ]r�4  (jw*  ]r�4  (jy*  ]r�4  (hh	e]r�4  (hh	e]r�4  (hjN  e]r�4  (j~*  ]r�4  (hh	e]r�4  (hhe]r�4  (hjN  e]r�4  (j�-  ]r�4  (hh	e]r�4  (hh	eeee]r�4  (hh&ee]r�4  (h]r�4  (hh e]r�4  (hhe]r�4  (hh	e]r�4  (h%heeej�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  ]r�4  (ju*  ]r�4  (jw*  ]r�4  (jy*  ]r�4  (hh	e]r�4  (hh	e]r�4  (hjN  e]r�4  (j~*  ]r�4  (hh	e]r�4  (hhe]r�4  (hjN  e]r�4  (j�-  ]r�4  (hh	e]r�4  (hh	eeee]r�4  (hh&ee]r�4  (h]r�4  (hh e]r�4  (hhe]r�4  (hh	e]r�4  (h%heeej�4  j�4  ]r�4  (ju*  ]r�4  (jw*  ]r�4  (jy*  ]r�4  (hh	e]r�4  (hh	e]r�4  (hjN  e]r�4  (j~*  ]r�4  (hh	e]r�4  (hhe]r�4  (hjN  e]r�4  (j�-  ]r�4  (hh	e]r�4  (hh	eeee]r�4  (hh&ee]r�4  (h]r�4  (hh e]r�4  (hhe]r�4  (hh	e]r�4  (h%heeej�4  j�4  j�4  ]r�4  (ju*  ]r�4  (jw*  ]r�4  (jy*  ]r�4  (hh	e]r�4  (hh	e]r�4  (hjN  e]r�4  (j~*  ]r�4  (hh	e]r�4  (hhe]r�4  (hjN  e]r�4  (j�-  ]r�4  (hh	e]r�4  (hh	eeee]r�4  (hh&ee]r�4  (h]r 5  (hh e]r5  (hhe]r5  (hh	e]r5  (h%heeej�4  j�4  ]r5  (ju*  ]r5  (jw*  ]r5  (jy*  ]r5  (hh	e]r5  (hh	e]r	5  (hjN  e]r
5  (j~*  ]r5  (hh	e]r5  (hhe]r5  (hjN  e]r5  (j�-  ]r5  (hh	e]r5  (hh	eeee]r5  (hh&ee]r5  (h]r5  (hh e]r5  (hhe]r5  (hh	e]r5  (h%heeej5  j5  j5  j5  ]r5  (ju*  ]r5  (jw*  ]r5  (jy*  ]r5  (hh	e]r5  (hh	e]r5  (hjN  e]r5  (j~*  ]r5  (hh	e]r5  (hhe]r 5  (hjN  e]r!5  (j�-  ]r"5  (hh	e]r#5  (hh	eeee]r$5  (hh&ee]r%5  (h]r&5  (hh e]r'5  (hhe]r(5  (hh	e]r)5  (h%heeej5  j5  ]r*5  (ju*  ]r+5  (jw*  ]r,5  (jy*  ]r-5  (hh	e]r.5  (hh	e]r/5  (hjN  e]r05  (j~*  ]r15  (hh	e]r25  (hhe]r35  (hjN  e]r45  (j�-  ]r55  (hh	e]r65  (hh	eeee]r75  (hh&ee]r85  (h]r95  (hh e]r:5  (hhe]r;5  (hh	e]r<5  (h%heeej*5  j*5  j*5  j*5  j*5  j*5  j*5  j*5  ]r=5  (ju*  ]r>5  (jw*  ]r?5  (jy*  ]r@5  (hh	e]rA5  (hh	e]rB5  (hjN  e]rC5  (j~*  ]rD5  (hh	e]rE5  (hhe]rF5  (hjN  e]rG5  (j�-  ]rH5  (hh	e]rI5  (hh	eeee]rJ5  (hh&ee]rK5  (h]rL5  (hh e]rM5  (hhe]rN5  (hh	e]rO5  (h%heeej=5  ]rP5  (ju*  ]rQ5  (jw*  ]rR5  (jy*  ]rS5  (hh	e]rT5  (hh	e]rU5  (hjN  e]rV5  (j~*  ]rW5  (hh	e]rX5  (hhe]rY5  (hjN  e]rZ5  (j�-  ]r[5  (hh	e]r\5  (hh	eeee]r]5  (hh&ee]r^5  (h]r_5  (hh e]r`5  (hhe]ra5  (hh	e]rb5  (h%heee]rc5  (ju*  ]rd5  (jw*  ]re5  (jy*  ]rf5  (hh	e]rg5  (hh	e]rh5  (hjN  e]ri5  (j~*  ]rj5  (hh	e]rk5  (hhe]rl5  (hjN  e]rm5  (j�-  ]rn5  (hh	e]ro5  (hh	eeee]rp5  (hh&ee]rq5  (h]rr5  (hh e]rs5  (hhe]rt5  (hh	e]ru5  (h%heee]rv5  (ju*  ]rw5  (jw*  ]rx5  (jy*  ]ry5  (hh	e]rz5  (hh	e]r{5  (hjN  e]r|5  (j~*  ]r}5  (hh	e]r~5  (hhe]r5  (hjN  e]r�5  (j�-  ]r�5  (hh	e]r�5  (hh	eeee]r�5  (hh&ee]r�5  (h]r�5  (hh e]r�5  (hhe]r�5  (hh	e]r�5  (h%heee]r�5  (ju*  ]r�5  (jw*  ]r�5  (jy*  ]r�5  (hh	e]r�5  (hh	e]r�5  (hjN  e]r�5  (j~*  ]r�5  (hh	e]r�5  (hhe]r�5  (hjN  e]r�5  (j�-  ]r�5  (hh	e]r�5  (hh	eeee]r�5  (hh&ee]r�5  (h]r�5  (hh e]r�5  (hhe]r�5  (hh	e]r�5  (h%heee]r�5  (ju*  ]r�5  (jw*  ]r�5  (jy*  ]r�5  (hh	e]r�5  (hh	e]r�5  (hjN  e]r�5  (j~*  ]r�5  (hh	e]r�5  (hhe]r�5  (hjN  e]r�5  (j�-  ]r�5  (hh	e]r�5  (hh	eeee]r�5  (hh&ee]r�5  (h]r�5  (hh e]r�5  (hhe]r�5  (hh	e]r�5  (h%heee]r�5  (ju*  ]r�5  (jw*  ]r�5  (jy*  ]r�5  (hh	e]r�5  (hh	e]r�5  (hjN  e]r�5  (j~*  ]r�5  (hhe]r�5  (hhe]r�5  (hjN  e]r�5  (j�-  ]r�5  (hh	e]r�5  (hh	eeee]r�5  (hh&ee]r�5  (h]r�5  (hh e]r�5  (hhe]r�5  (hh	e]r�5  (h%heeej�5  j�5  j�5  j�5  j�5  ]r�5  (ju*  ]r�5  (jw*  ]r�5  (jy*  ]r�5  (hh	e]r�5  (hh	e]r�5  (hjN  e]r�5  (j~*  ]r�5  (hhe]r�5  (hhe]r�5  (hjN  e]r�5  (j�-  ]r�5  (hh	e]r�5  (hh	eeee]r�5  (hh&ee]r�5  (h]r�5  (hh e]r�5  (hhe]r�5  (hhe]r�5  (h%heee]r�5  (ju*  ]r�5  (jw*  ]r�5  (jy*  ]r�5  (hh	e]r�5  (hh	e]r�5  (hjN  e]r�5  (j~*  ]r�5  (hhe]r�5  (hhe]r�5  (hjN  e]r�5  (j�-  ]r�5  (hh	e]r�5  (hh	eeee]r�5  (hh&ee]r�5  (h]r�5  (hh e]r�5  (hhe]r�5  (hh	e]r�5  (h%heee]r�5  (ju*  ]r�5  (jw*  ]r�5  (jy*  ]r�5  (hh	e]r�5  (hh	e]r�5  (hjN  e]r�5  (j~*  ]r�5  (hh	e]r�5  (hhe]r�5  (hjN  e]r�5  (j�-  ]r�5  (hh	e]r�5  (hh	eeee]r�5  (hh&ee]r�5  (h]r�5  (hh e]r�5  (hhe]r�5  (hh	e]r�5  (h%heeej�5  j�5  j�5  j�5  j�5  ]r�5  (ju*  ]r�5  (jw*  ]r�5  (jy*  ]r�5  (hh	e]r�5  (hh	e]r 6  (hjN  e]r6  (j~*  ]r6  (hh	e]r6  (hhe]r6  (hjN  e]r6  (j�-  ]r6  (hh	e]r6  (hh	eeee]r6  (hh&ee]r	6  (h]r
6  (hh e]r6  (hhe]r6  (hh	e]r6  (h%heeej�5  ]r6  (ju*  ]r6  (jw*  ]r6  (jy*  ]r6  (hh	e]r6  (hh	e]r6  (hjN  e]r6  (j~*  ]r6  (hh	e]r6  (hhe]r6  (hjN  e]r6  (j�-  ]r6  (hh	e]r6  (hh	eeee]r6  (hh&ee]r6  (h]r6  (hh e]r6  (hhe]r6  (hh	e]r 6  (h%heee]r!6  (ju*  ]r"6  (jw*  ]r#6  (jy*  ]r$6  (hh	e]r%6  (hh	e]r&6  (hjN  e]r'6  (j~*  ]r(6  (hh	e]r)6  (hhe]r*6  (hjN  e]r+6  (j�-  ]r,6  (hh	e]r-6  (hh	eeee]r.6  (hh&ee]r/6  (h]r06  (hh e]r16  (hhe]r26  (hh	e]r36  (h%heeej!6  j!6  j!6  j!6  ]r46  (ju*  ]r56  (jw*  ]r66  (jy*  ]r76  (hh	e]r86  (hh	e]r96  (hjN  e]r:6  (j~*  ]r;6  (hh	e]r<6  (hhe]r=6  (hjN  e]r>6  (j�-  ]r?6  (hh	e]r@6  (hh	eeee]rA6  (hh&ee]rB6  (h]rC6  (hh e]rD6  (hhe]rE6  (hh	e]rF6  (h%heee]rG6  (ju*  ]rH6  (jw*  ]rI6  (jy*  ]rJ6  (hh	e]rK6  (hh	e]rL6  (hjN  e]rM6  (j~*  ]rN6  (hh	e]rO6  (hhe]rP6  (hjN  e]rQ6  (j�-  ]rR6  (hh	e]rS6  (hh	eeee]rT6  (hh&ee]rU6  (h]rV6  (hh e]rW6  (hhe]rX6  (hh	e]rY6  (h%heeejG6  ]rZ6  (ju*  ]r[6  (jw*  ]r\6  (jy*  ]r]6  (hh	e]r^6  (hh	e]r_6  (hjN  e]r`6  (j~*  ]ra6  (hh	e]rb6  (hhe]rc6  (hjN  e]rd6  (j�-  ]re6  (hh	e]rf6  (hh	eeee]rg6  (hh&ee]rh6  (h]ri6  (hh e]rj6  (hhe]rk6  (hh	e]rl6  (h%heeejZ6  jZ6  jZ6  jZ6  jZ6  ]rm6  (ju*  ]rn6  (jw*  ]ro6  (jy*  ]rp6  (hh	e]rq6  (hh	e]rr6  (hjN  e]rs6  (j~*  ]rt6  (hh	e]ru6  (hhe]rv6  (hjN  e]rw6  (j�-  ]rx6  (hh	e]ry6  (hh	eeee]rz6  (hh&ee]r{6  (h]r|6  (hh e]r}6  (hhe]r~6  (hh	e]r6  (h%heeejm6  jm6  jm6  ]r�6  (ju*  ]r�6  (jw*  ]r�6  (jy*  ]r�6  (hh	e]r�6  (hh	e]r�6  (hjN  e]r�6  (j~*  ]r�6  (hh	e]r�6  (hhe]r�6  (hjN  e]r�6  (j�-  ]r�6  (hh	e]r�6  (hh	eeee]r�6  (hh&ee]r�6  (h]r�6  (hh e]r�6  (hhe]r�6  (hh	e]r�6  (h%heeej�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  ]r�6  (ju*  ]r�6  (jw*  ]r�6  (jy*  ]r�6  (hh	e]r�6  (hh	e]r�6  (hjN  e]r�6  (j~*  ]r�6  (hh	e]r�6  (hhe]r�6  (hjN  e]r�6  (j�-  ]r�6  (hh	e]r�6  (hh	eeee]r�6  (hh&ee]r�6  (h]r�6  (hh e]r�6  (hhe]r�6  (hh	e]r�6  (h%heee]r�6  (ju*  ]r�6  (jw*  ]r�6  (jy*  ]r�6  (hh	e]r�6  (hh	e]r�6  (hjN  e]r�6  (j~*  ]r�6  (hh	e]r�6  (hhe]r�6  (hjN  e]r�6  (j�-  ]r�6  (hh	e]r�6  (hh	eeee]r�6  (hh&ee]r�6  (h]r�6  (hh e]r�6  (hhe]r�6  (hh	e]r�6  (h%heeej�6  j�6  j�6  ]r�6  (ju*  ]r�6  (jw*  ]r�6  (jy*  ]r�6  (hh	e]r�6  (hh	e]r�6  (hjN  e]r�6  (j~*  ]r�6  (hh	e]r�6  (hhe]r�6  (hjN  e]r�6  (j�-  ]r�6  (hh	e]r�6  (hh	eeee]r�6  (hh&ee]r�6  (h]r�6  (hh e]r�6  (hhe]r�6  (hh	e]r�6  (h%heee]r�6  (ju*  ]r�6  (jw*  ]r�6  (jy*  ]r�6  (hh	e]r�6  (hh	e]r�6  (hjN  e]r�6  (j~*  ]r�6  (hh	e]r�6  (hhe]r�6  (hjN  e]r�6  (j�-  ]r�6  (hh	e]r�6  (hh	eeee]r�6  (hh&ee]r�6  (h]r�6  (hh e]r�6  (hhe]r�6  (hh	e]r�6  (h%heeej�6  ]r�6  (ju*  ]r�6  (jw*  ]r�6  (jy*  ]r�6  (hh	e]r�6  (hh	e]r�6  (hjN  e]r�6  (j~*  ]r�6  (hhe]r�6  (hhe]r�6  (hjN  e]r�6  (j�-  ]r�6  (hh	e]r�6  (hh	eeee]r�6  (hh&ee]r�6  (h]r�6  (hh e]r�6  (hhe]r�6  (hh	e]r�6  (h%heeej�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  ]r�6  (ju*  ]r�6  (jw*  ]r�6  (jy*  ]r�6  (hh	e]r�6  (hh	e]r�6  (hjN  e]r�6  (j~*  ]r�6  (hhe]r�6  (hhe]r�6  (hjN  e]r�6  (j�-  ]r�6  (hh	e]r�6  (hh	eeee]r�6  (hh&ee]r 7  (h]r7  (hh e]r7  (hhe]r7  (hh	e]r7  (h%heeej�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  ]r7  (ju*  ]r7  (jw*  ]r7  (jy*  ]r7  (hh	e]r	7  (hh	e]r
7  (hjN  e]r7  (j~*  ]r7  (hhe]r7  (hhe]r7  (hjN  e]r7  (j�-  ]r7  (hh	e]r7  (hh	eeee]r7  (hh&ee]r7  (h]r7  (hh e]r7  (hhe]r7  (hh	e]r7  (h%heeej7  j7  j7  j7  j7  ]r7  (ju*  ]r7  (jw*  ]r7  (jy*  ]r7  (hh	e]r7  (hh	e]r7  (hjN  e]r7  (j~*  ]r7  (hhe]r 7  (hhe]r!7  (hjN  e]r"7  (j�-  ]r#7  (hh	e]r$7  (hh	eeee]r%7  (hh&ee]r&7  (h]r'7  (hh e]r(7  (hhe]r)7  (hh	e]r*7  (h%heeej7  j7  j7  j7  ]r+7  (ju*  ]r,7  (jw*  ]r-7  (jy*  ]r.7  (hh	e]r/7  (hh	e]r07  (hjN  e]r17  (j~*  ]r27  (hhe]r37  (hhe]r47  (hjN  e]r57  (j�-  ]r67  (hh	e]r77  (hh	eeee]r87  (hh&ee]r97  (h]r:7  (hh e]r;7  (hhe]r<7  (hh	e]r=7  (h%heeej+7  j+7  j+7  ]r>7  (ju*  ]r?7  (jw*  ]r@7  (jy*  ]rA7  (hh	e]rB7  (hh	e]rC7  (hjN  e]rD7  (j~*  ]rE7  (hhe]rF7  (hhe]rG7  (hjN  e]rH7  (j�-  ]rI7  (hh	e]rJ7  (hh	eeee]rK7  (hh&ee]rL7  (h]rM7  (hh e]rN7  (hhe]rO7  (hh	e]rP7  (h%heeej>7  j>7  j>7  j>7  j>7  ]rQ7  (ju*  ]rR7  (jw*  ]rS7  (jy*  ]rT7  (hh	e]rU7  (hh	e]rV7  (hjN  e]rW7  (j~*  ]rX7  (hhe]rY7  (hhe]rZ7  (hjN  e]r[7  (j�-  ]r\7  (hh	e]r]7  (hh	eeee]r^7  (hh&ee]r_7  (h]r`7  (hh e]ra7  (hhe]rb7  (hh	e]rc7  (h%heeejQ7  jQ7  jQ7  jQ7  jQ7  jQ7  jQ7  jQ7  ]rd7  (ju*  ]re7  (jw*  ]rf7  (jy*  ]rg7  (hh	e]rh7  (hh	e]ri7  (hjN  e]rj7  (j~*  ]rk7  (hhe]rl7  (hhe]rm7  (hjN  e]rn7  (j�-  ]ro7  (hh	e]rp7  (hh	eeee]rq7  (hh&ee]rr7  (h]rs7  (hh e]rt7  (hhe]ru7  (hh	e]rv7  (h%heeejd7  jd7  jd7  jd7  jd7  ]rw7  (ju*  ]rx7  (jw*  ]ry7  (jy*  ]rz7  (hh	e]r{7  (hh	e]r|7  (hjN  e]r}7  (j~*  ]r~7  (hhe]r7  (hhe]r�7  (hjN  e]r�7  (j�-  ]r�7  (hh	e]r�7  (hh	eeee]r�7  (hh&ee]r�7  (h]r�7  (hh e]r�7  (hhe]r�7  (hh	e]r�7  (h%heeejw7  jw7  jw7  jw7  jw7  jw7  jw7  jw7  jw7  jw7  ]r�7  (ju*  ]r�7  (jw*  ]r�7  (jy*  ]r�7  (hh	e]r�7  (hh	e]r�7  (hjN  e]r�7  (j~*  ]r�7  (hhe]r�7  (hhe]r�7  (hjN  e]r�7  (j�-  ]r�7  (hh	e]r�7  (hh	eeee]r�7  (hh&ee]r�7  (h]r�7  (hh e]r�7  (hhe]r�7  (hh	e]r�7  (h%heeej�7  ]r�7  (ju*  ]r�7  (jw*  ]r�7  (jy*  ]r�7  (hh	e]r�7  (hh	e]r�7  (hjN  e]r�7  (j~*  ]r�7  (hhe]r�7  (hhe]r�7  (hjN  e]r�7  (j�-  ]r�7  (hh	e]r�7  (hh	eeee]r�7  (hh&ee]r�7  (h]r�7  (hh e]r�7  (hhe]r�7  (hh	e]r�7  (h%heee]r�7  (ju*  ]r�7  (jw*  ]r�7  (jy*  ]r�7  (hh	e]r�7  (hh	e]r�7  (hjN  e]r�7  (j~*  ]r�7  (hhe]r�7  (hhe]r�7  (hjN  e]r�7  (j�-  ]r�7  (hh	e]r�7  (hh	eeee]r�7  (hh&ee]r�7  (h]r�7  (hh e]r�7  (hhe]r�7  (hh	e]r�7  (h%heee]r�7  (ju*  ]r�7  (jw*  ]r�7  (jy*  ]r�7  (hh	e]r�7  (hh	e]r�7  (hjN  e]r�7  (j~*  ]r�7  (hhe]r�7  (hhe]r�7  (hjN  e]r�7  (j�-  ]r�7  (hh	e]r�7  (hh	eeee]r�7  (hh&ee]r�7  (h]r�7  (hh e]r�7  (hhe]r�7  (hh	e]r�7  (h%heeej�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  ]r�7  (ju*  ]r�7  (jw*  ]r�7  (jy*  ]r�7  (hh	e]r�7  (hh	e]r�7  (hjN  e]r�7  (j~*  ]r�7  (hhe]r�7  (hhe]r�7  (hjN  e]r�7  (j�-  ]r�7  (hh	e]r�7  (hh	eeee]r�7  (hh&ee]r�7  (h]r�7  (hh e]r�7  (hhe]r�7  (hh	e]r�7  (h%heeej�7  j�7  j�7  j�7  j�7  ]r�7  (ju*  ]r�7  (jw*  ]r�7  (jy*  ]r�7  (hh	e]r�7  (hh	e]r�7  (hjN  e]r�7  (j~*  ]r�7  (hhe]r�7  (hhe]r�7  (hjN  e]r�7  (j�-  ]r�7  (hh	e]r�7  (hh	eeee]r�7  (hh&ee]r�7  (h]r�7  (hh e]r�7  (hhe]r�7  (hh	e]r�7  (h%heeej�7  j�7  ]r�7  (ju*  ]r�7  (jw*  ]r�7  (jy*  ]r�7  (hh	e]r 8  (hh	e]r8  (hjN  e]r8  (j~*  ]r8  (hhe]r8  (hhe]r8  (hjN  e]r8  (j�-  ]r8  (hh	e]r8  (hh	eeee]r	8  (hh&ee]r
8  (h]r8  (hh e]r8  (hhe]r8  (hh	e]r8  (h%heee]r8  (ju*  ]r8  (jw*  ]r8  (jy*  ]r8  (hh	e]r8  (hh	e]r8  (hjN  e]r8  (j~*  ]r8  (hhe]r8  (hhe]r8  (hjN  e]r8  (j�-  ]r8  (hh	e]r8  (hh	eeee]r8  (hh&ee]r8  (h]r8  (hh e]r8  (hhe]r 8  (hh	e]r!8  (h%heee]r"8  (ju*  ]r#8  (jw*  ]r$8  (jy*  ]r%8  (hh	e]r&8  (hh	e]r'8  (hjN  e]r(8  (j~*  ]r)8  (hhe]r*8  (hhe]r+8  (hjN  e]r,8  (j�-  ]r-8  (hh	e]r.8  (hh	eeee]r/8  (hh&ee]r08  (h]r18  (hh e]r28  (hhe]r38  (hh	e]r48  (h%heee]r58  (ju*  ]r68  (jw*  ]r78  (jy*  ]r88  (hh	e]r98  (hh	e]r:8  (hjN  e]r;8  (j~*  ]r<8  (hhe]r=8  (hhe]r>8  (hjN  e]r?8  (j�-  ]r@8  (hh	e]rA8  (hh	eeee]rB8  (hh&ee]rC8  (h]rD8  (hh e]rE8  (hhe]rF8  (hh	e]rG8  (h%heee]rH8  (ju*  ]rI8  (jw*  ]rJ8  (jy*  ]rK8  (hh	e]rL8  (hh	e]rM8  (hjN  e]rN8  (j~*  ]rO8  (hhe]rP8  (hhe]rQ8  (hjN  e]rR8  (j�-  ]rS8  (hh	e]rT8  (hh	eeee]rU8  (hh&ee]rV8  (h]rW8  (hh e]rX8  (hhe]rY8  (hh	e]rZ8  (h%heeejH8  jH8  jH8  ]r[8  (ju*  ]r\8  (jw*  ]r]8  (jy*  ]r^8  (hh	e]r_8  (hh	e]r`8  (hjN  e]ra8  (j~*  ]rb8  (hhe]rc8  (hhe]rd8  (hjN  e]re8  (j�-  ]rf8  (hh	e]rg8  (hh	eeee]rh8  (hh&ee]ri8  (h]rj8  (hh e]rk8  (hhe]rl8  (hh	e]rm8  (h%heeej[8  j[8  j[8  j[8  j[8  j[8  ]rn8  (ju*  ]ro8  (jw*  ]rp8  (jy*  ]rq8  (hh	e]rr8  (hh	e]rs8  (hjN  e]rt8  (j~*  ]ru8  (hhe]rv8  (hhe]rw8  (hjN  e]rx8  (j�-  ]ry8  (hh	e]rz8  (hh	eeee]r{8  (hh&ee]r|8  (h]r}8  (hh e]r~8  (hhe]r8  (hh	e]r�8  (h%heee]r�8  (ju*  ]r�8  (jw*  ]r�8  (jy*  ]r�8  (hh	e]r�8  (hh	e]r�8  (hjN  e]r�8  (j~*  ]r�8  (hhe]r�8  (hhe]r�8  (hjN  e]r�8  (j�-  ]r�8  (hh	e]r�8  (hh	eeee]r�8  (hh&ee]r�8  (h]r�8  (hh e]r�8  (hhe]r�8  (hh	e]r�8  (h%heeej�8  j�8  ]r�8  (ju*  ]r�8  (jw*  ]r�8  (jy*  ]r�8  (hh	e]r�8  (hh	e]r�8  (hjN  e]r�8  (j~*  ]r�8  (hhe]r�8  (hhe]r�8  (hjN  e]r�8  (j�-  ]r�8  (hh	e]r�8  (hh	eeee]r�8  (hh&ee]r�8  (h]r�8  (hh e]r�8  (hhe]r�8  (hh	e]r�8  (h%heeej�8  ]r�8  (ju*  ]r�8  (jw*  ]r�8  (jy*  ]r�8  (hh	e]r�8  (hh	e]r�8  (hjN  e]r�8  (j~*  ]r�8  (hhe]r�8  (hhe]r�8  (hjN  e]r�8  (j�-  ]r�8  (hh	e]r�8  (hh	eeee]r�8  (hh&ee]r�8  (h]r�8  (hh e]r�8  (hhe]r�8  (hh	e]r�8  (h%heee]r�8  (ju*  ]r�8  (jw*  ]r�8  (jy*  ]r�8  (hh	e]r�8  (hh	e]r�8  (hjN  e]r�8  (j~*  ]r�8  (hhe]r�8  (hhe]r�8  (hjN  e]r�8  (j�-  ]r�8  (hh	e]r�8  (hh	eeee]r�8  (hh&ee]r�8  (h]r�8  (hh e]r�8  (hhe]r�8  (hhe]r�8  (h%heeej�8  j�8  j�8  j�8  j�8  j�8  ]r�8  (ju*  ]r�8  (jw*  ]r�8  (jy*  ]r�8  (hh	e]r�8  (hh	e]r�8  (hjN  e]r�8  (j~*  ]r�8  (hhe]r�8  (hhe]r�8  (hjN  e]r�8  (j�-  ]r�8  (hh	e]r�8  (hh	eeee]r�8  (hh&ee]r�8  (h]r�8  (hh e]r�8  (hhe]r�8  (hhe]r�8  (h%heeej�8  j�8  ]r�8  (ju*  ]r�8  (jw*  ]r�8  (jy*  ]r�8  (hh	e]r�8  (hh	e]r�8  (hjN  e]r�8  (j~*  ]r�8  (hhe]r�8  (hhe]r�8  (hjN  e]r�8  (j�-  ]r�8  (hh	e]r�8  (hh	eeee]r�8  (hh&ee]r�8  (h]r�8  (hh e]r�8  (hhe]r�8  (hhe]r�8  (h%heeej�8  j�8  j�8  j�8  j�8  j�8  j�8  j�8  j�8  ]r�8  (ju*  ]r�8  (jw*  ]r�8  (jy*  ]r�8  (hh	e]r�8  (hh	e]r�8  (hjN  e]r�8  (j~*  ]r�8  (hhe]r�8  (hhe]r�8  (hjN  e]r�8  (j�-  ]r�8  (hh	e]r�8  (hh	eeee]r 9  (hh&ee]r9  (h]r9  (hh e]r9  (hhe]r9  (hhe]r9  (h%heeej�8  j�8  j�8  ]r9  (ju*  ]r9  (jw*  ]r9  (jy*  ]r	9  (hh	e]r
9  (hh	e]r9  (hjN  e]r9  (j~*  ]r9  (hh	e]r9  (hhe]r9  (hjN  e]r9  (j�-  ]r9  (hh	e]r9  (hh	eeee]r9  (hh&ee]r9  (h]r9  (hh e]r9  (hhe]r9  (hhe]r9  (h%heeej9  ]r9  (ju*  ]r9  (jw*  ]r9  (jy*  ]r9  (hh	e]r9  (hh	e]r9  (hjN  e]r9  (j~*  ]r 9  (hh	e]r!9  (hhe]r"9  (hjN  e]r#9  (j�-  ]r$9  (hh	e]r%9  (hh	eeee]r&9  (hh&ee]r'9  (h]r(9  (hh e]r)9  (hhe]r*9  (hhe]r+9  (h%heeej9  j9  j9  j9  j9  ]r,9  (ju*  ]r-9  (jw*  ]r.9  (jy*  ]r/9  (hh	e]r09  (hh	e]r19  (hjN  e]r29  (j~*  ]r39  (hh	e]r49  (hhe]r59  (hjN  e]r69  (j�-  ]r79  (hh	e]r89  (hh	eeee]r99  (hh&ee]r:9  (h]r;9  (hh e]r<9  (hhe]r=9  (hhe]r>9  (h%heeej,9  j,9  j,9  j,9  ]r?9  (ju*  ]r@9  (jw*  ]rA9  (jy*  ]rB9  (hh	e]rC9  (hh	e]rD9  (hjN  e]rE9  (j~*  ]rF9  (hh	e]rG9  (hhe]rH9  (hjN  e]rI9  (j�-  ]rJ9  (hh	e]rK9  (hh	eeee]rL9  (hh&ee]rM9  (h]rN9  (hh e]rO9  (hhe]rP9  (hhe]rQ9  (h%heee]rR9  (ju*  ]rS9  (jw*  ]rT9  (jy*  ]rU9  (hh	e]rV9  (hh	e]rW9  (hjN  e]rX9  (j~*  ]rY9  (hh	e]rZ9  (hhe]r[9  (hjN  e]r\9  (j�-  ]r]9  (hh	e]r^9  (hh	eeee]r_9  (hh&ee]r`9  (h]ra9  (hh e]rb9  (hhe]rc9  (hhe]rd9  (h%heeejR9  jR9  jR9  jR9  jR9  jR9  jR9  jR9  ]re9  (ju*  ]rf9  (jw*  ]rg9  (jy*  ]rh9  (hh	e]ri9  (hh	e]rj9  (hjN  e]rk9  (j~*  ]rl9  (hh	e]rm9  (hhe]rn9  (hjN  e]ro9  (j�-  ]rp9  (hh	e]rq9  (hh	eeee]rr9  (hh&ee]rs9  (h]rt9  (hh e]ru9  (hhe]rv9  (hh	e]rw9  (h%heeeje9  je9  je9  je9  je9  je9  je9  je9  je9  je9  ]rx9  (ju*  ]ry9  (jw*  ]rz9  (jy*  ]r{9  (hh	e]r|9  (hh	e]r}9  (hjN  e]r~9  (j~*  ]r9  (hh	e]r�9  (hhe]r�9  (hjN  e]r�9  (j�-  ]r�9  (hh	e]r�9  (hh	eeee]r�9  (hh&ee]r�9  (h]r�9  (hh e]r�9  (hhe]r�9  (hh	e]r�9  (h%heee]r�9  (ju*  ]r�9  (jw*  ]r�9  (jy*  ]r�9  (hh	e]r�9  (hh	e]r�9  (hjN  e]r�9  (j~*  ]r�9  (hh	e]r�9  (hhe]r�9  (hjN  e]r�9  (j�-  ]r�9  (hh	e]r�9  (hh	eeee]r�9  (hh&ee]r�9  (h]r�9  (hh e]r�9  (hhe]r�9  (hh	e]r�9  (h%heeej�9  j�9  ]r�9  (ju*  ]r�9  (jw*  ]r�9  (jy*  ]r�9  (hh	e]r�9  (hh	e]r�9  (hjN  e]r�9  (j~*  ]r�9  (hh	e]r�9  (hhe]r�9  (hjN  e]r�9  (j�-  ]r�9  (hh	e]r�9  (hh	eeee]r�9  (hh&ee]r�9  (h]r�9  (hh e]r�9  (hhe]r�9  (hh	e]r�9  (h%heee]r�9  (ju*  ]r�9  (jw*  ]r�9  (jy*  ]r�9  (hh	e]r�9  (hh	e]r�9  (hjN  e]r�9  (j~*  ]r�9  (hhe]r�9  (hhe]r�9  (hjN  e]r�9  (j�-  ]r�9  (hh	e]r�9  (hh	eeee]r�9  (hh&ee]r�9  (h]r�9  (hh e]r�9  (hhe]r�9  (hh	e]r�9  (h%heeej�9  j�9  ]r�9  (ju*  ]r�9  (jw*  ]r�9  (jy*  ]r�9  (hh	e]r�9  (hh	e]r�9  (hjN  e]r�9  (j~*  ]r�9  (hhe]r�9  (hhe]r�9  (hjN  e]r�9  (j�-  ]r�9  (hh	e]r�9  (hh	eeee]r�9  (hh&ee]r�9  (h]r�9  (hh e]r�9  (hhe]r�9  (hh	e]r�9  (h%heeej�9  j�9  j�9  j�9  ]r�9  (ju*  ]r�9  (jw*  ]r�9  (jy*  ]r�9  (hh	e]r�9  (hh	e]r�9  (hjN  e]r�9  (j~*  ]r�9  (hhe]r�9  (hhe]r�9  (hjN  e]r�9  (j�-  ]r�9  (hh	e]r�9  (hh	eeee]r�9  (hh&ee]r�9  (h]r�9  (hh e]r�9  (hhe]r�9  (hh	e]r�9  (h%heeej�9  j�9  ]r�9  (ju*  ]r�9  (jw*  ]r�9  (jy*  ]r�9  (hh	e]r�9  (hh	e]r�9  (hjN  e]r�9  (j~*  ]r�9  (hhe]r�9  (hhe]r�9  (hjN  e]r�9  (j�-  ]r�9  (hh	e]r�9  (hh	eeee]r�9  (hh&ee]r�9  (h]r�9  (hh e]r�9  (hhe]r�9  (hh	e]r�9  (h%heee]r�9  (ju*  ]r�9  (jw*  ]r�9  (jy*  ]r :  (hh	e]r:  (hh	e]r:  (hjN  e]r:  (j~*  ]r:  (hhe]r:  (hhe]r:  (hjN  e]r:  (j�-  ]r:  (hh	e]r	:  (hh	eeee]r
:  (hh&ee]r:  (h]r:  (hh e]r:  (hhe]r:  (hh	e]r:  (h%heeej�9  j�9  j�9  j�9  j�9  ]r:  (ju*  ]r:  (jw*  ]r:  (jy*  ]r:  (hh	e]r:  (hh	e]r:  (hjN  e]r:  (j~*  ]r:  (hhe]r:  (hhe]r:  (hjN  e]r:  (j�-  ]r:  (hh	e]r:  (hh	eeee]r:  (hh&ee]r:  (h]r:  (hh e]r :  (hhe]r!:  (hh	e]r":  (h%heeej:  j:  j:  j:  j:  j:  ]r#:  (ju*  ]r$:  (jw*  ]r%:  (jy*  ]r&:  (hh	e]r':  (hh	e]r(:  (hjN  e]r):  (j~*  ]r*:  (hhe]r+:  (hhe]r,:  (hjN  e]r-:  (j�-  ]r.:  (hh	e]r/:  (hh	eeee]r0:  (hh&ee]r1:  (h]r2:  (hh e]r3:  (hhe]r4:  (hh	e]r5:  (h%heeej#:  j#:  j#:  ]r6:  (ju*  ]r7:  (jw*  ]r8:  (jy*  ]r9:  (hh	e]r::  (hh	e]r;:  (hjN  e]r<:  (j~*  ]r=:  (hhe]r>:  (hhe]r?:  (hjN  e]r@:  (j�-  ]rA:  (hh	e]rB:  (hh	eeee]rC:  (hh&ee]rD:  (h]rE:  (hh e]rF:  (hhe]rG:  (hh	e]rH:  (h%heeej6:  j6:  j6:  ]rI:  (ju*  ]rJ:  (jw*  ]rK:  (jy*  ]rL:  (hh	e]rM:  (hh	e]rN:  (hjN  e]rO:  (j~*  ]rP:  (hhe]rQ:  (hhe]rR:  (hjN  e]rS:  (j�-  ]rT:  (hh	e]rU:  (hh	eeee]rV:  (hh&ee]rW:  (h]rX:  (hh e]rY:  (hhe]rZ:  (hh	e]r[:  (h%heee]r\:  (ju*  ]r]:  (jw*  ]r^:  (jy*  ]r_:  (hh	e]r`:  (hh	e]ra:  (hjN  e]rb:  (j~*  ]rc:  (hhe]rd:  (hhe]re:  (hjN  e]rf:  (j�-  ]rg:  (hh	e]rh:  (hh	eeee]ri:  (hh&ee]rj:  (h]rk:  (hh e]rl:  (hhe]rm:  (hh	e]rn:  (h%heeej\:  j\:  ]ro:  (ju*  ]rp:  (jw*  ]rq:  (jy*  ]rr:  (hh	e]rs:  (hh	e]rt:  (hjN  e]ru:  (j~*  ]rv:  (hhe]rw:  (hhe]rx:  (hjN  e]ry:  (j�-  ]rz:  (hh	e]r{:  (hh	eeee]r|:  (hh&ee]r}:  (h]r~:  (hh e]r:  (hhe]r�:  (hh	e]r�:  (h%heeejo:  jo:  jo:  ]r�:  (ju*  ]r�:  (jw*  ]r�:  (jy*  ]r�:  (hh	e]r�:  (hh	e]r�:  (hjN  e]r�:  (j~*  ]r�:  (hhe]r�:  (hhe]r�:  (hjN  e]r�:  (j�-  ]r�:  (hh	e]r�:  (hh	eeee]r�:  (hh&ee]r�:  (h]r�:  (hh e]r�:  (hhe]r�:  (hh	e]r�:  (h%heeej�:  ]r�:  (ju*  ]r�:  (jw*  ]r�:  (jy*  ]r�:  (hh	e]r�:  (hh	e]r�:  (hjN  e]r�:  (j~*  ]r�:  (hhe]r�:  (hhe]r�:  (hjN  e]r�:  (j�-  ]r�:  (hh	e]r�:  (hh	eeee]r�:  (hh&ee]r�:  (h]r�:  (hh e]r�:  (hhe]r�:  (hh	e]r�:  (h%heeej�:  j�:  j�:  ]r�:  (ju*  ]r�:  (jw*  ]r�:  (jy*  ]r�:  (hh	e]r�:  (hh	e]r�:  (hjN  e]r�:  (j~*  ]r�:  (hhe]r�:  (hhe]r�:  (hjN  e]r�:  (j�-  ]r�:  (hh	e]r�:  (hh	eeee]r�:  (hh&ee]r�:  (h]r�:  (hh e]r�:  (hhe]r�:  (hh	e]r�:  (h%heeej�:  j�:  j�:  ]r�:  (ju*  ]r�:  (jw*  ]r�:  (jy*  ]r�:  (hh	e]r�:  (hh	e]r�:  (hjN  e]r�:  (j~*  ]r�:  (hhe]r�:  (hhe]r�:  (hjN  e]r�:  (j�-  ]r�:  (hh	e]r�:  (hh	eeee]r�:  (hh&ee]r�:  (h]r�:  (hh e]r�:  (hhe]r�:  (hh	e]r�:  (h%heeej�:  j�:  ]r�:  (ju*  ]r�:  (jw*  ]r�:  (jy*  ]r�:  (hh	e]r�:  (hh	e]r�:  (hjN  e]r�:  (j~*  ]r�:  (hhe]r�:  (hhe]r�:  (hjN  e]r�:  (j�-  ]r�:  (hh	e]r�:  (hh	eeee]r�:  (hh&ee]r�:  (h]r�:  (hh e]r�:  (hhe]r�:  (hh	e]r�:  (h%heeej�:  j�:  j�:  j�:  j�:  j�:  ]r�:  (ju*  ]r�:  (jw*  ]r�:  (jy*  ]r�:  (hh	e]r�:  (hh	e]r�:  (hjN  e]r�:  (j~*  ]r�:  (hhe]r�:  (hhe]r�:  (hjN  e]r�:  (j�-  ]r�:  (hh	e]r�:  (hh	eeee]r�:  (hh&ee]r�:  (h]r�:  (hh e]r�:  (hhe]r�:  (hh	e]r�:  (h%heeej�:  j�:  ]r�:  (ju*  ]r�:  (jw*  ]r�:  (jy*  ]r�:  (hh	e]r�:  (hh	e]r�:  (hjN  e]r�:  (j~*  ]r�:  (hhe]r�:  (hhe]r�:  (hjN  e]r�:  (j�-  ]r�:  (hh	e]r ;  (hh	eeee]r;  (hh&ee]r;  (h]r;  (hh e]r;  (hhe]r;  (hh	e]r;  (h%heee]r;  (ju*  ]r;  (jw*  ]r	;  (jy*  ]r
;  (hh	e]r;  (hh	e]r;  (hjN  e]r;  (j~*  ]r;  (hhe]r;  (hhe]r;  (hjN  e]r;  (j�-  ]r;  (hh	e]r;  (hh	eeee]r;  (hh&ee]r;  (h]r;  (hh e]r;  (hhe]r;  (hhe]r;  (h%heeej;  j;  j;  j;  j;  j;  j;  j;  j;  j;  j;  ]r;  (ju*  ]r;  (jw*  ]r;  (jy*  ]r;  (hh	e]r;  (hh	e]r;  (hjN  e]r ;  (j~*  ]r!;  (hhe]r";  (hhe]r#;  (hjN  e]r$;  (j�-  ]r%;  (hh	e]r&;  (hh	eeee]r';  (hh&ee]r(;  (h]r);  (hh e]r*;  (hhe]r+;  (hhe]r,;  (h%heeej;  j;  j;  j;  j;  ]r-;  (ju*  ]r.;  (jw*  ]r/;  (jy*  ]r0;  (hh	e]r1;  (hh	e]r2;  (hjN  e]r3;  (j~*  ]r4;  (hhe]r5;  (hhe]r6;  (hjN  e]r7;  (j�-  ]r8;  (hh	e]r9;  (hh	eeee]r:;  (hh&ee]r;;  (h]r<;  (hh e]r=;  (hhe]r>;  (hhe]r?;  (h%heeej-;  j-;  j-;  ]r@;  (ju*  ]rA;  (jw*  ]rB;  (jy*  ]rC;  (hh	e]rD;  (hh	e]rE;  (hjN  e]rF;  (j~*  ]rG;  (hhe]rH;  (hhe]rI;  (hjN  e]rJ;  (j�-  ]rK;  (hh	e]rL;  (hh	eeee]rM;  (hh&ee]rN;  (h]rO;  (hh e]rP;  (hhe]rQ;  (hhe]rR;  (h%heeej@;  j@;  ]rS;  (ju*  ]rT;  (jw*  ]rU;  (jy*  ]rV;  (hh	e]rW;  (hh	e]rX;  (hjN  e]rY;  (j~*  ]rZ;  (hhe]r[;  (hhe]r\;  (hjN  e]r];  (j�-  ]r^;  (hh	e]r_;  (hh	eeee]r`;  (hh&ee]ra;  (h]rb;  (hh e]rc;  (hhe]rd;  (hh	e]re;  (h%heeejS;  jS;  ]rf;  (ju*  ]rg;  (jw*  ]rh;  (jy*  ]ri;  (hh	e]rj;  (hh	e]rk;  (hjN  e]rl;  (j~*  ]rm;  (hhe]rn;  (hhe]ro;  (hjN  e]rp;  (j�-  ]rq;  (hh	e]rr;  (hh	eeee]rs;  (hh&ee]rt;  (h]ru;  (hh e]rv;  (hhe]rw;  (hh	e]rx;  (h%heeejf;  jf;  ]ry;  (ju*  ]rz;  (jw*  ]r{;  (jy*  ]r|;  (hh	e]r};  (hh	e]r~;  (hjN  e]r;  (j~*  ]r�;  (hhe]r�;  (hhe]r�;  (hjN  e]r�;  (j�-  ]r�;  (hh	e]r�;  (hh	eeee]r�;  (hh&ee]r�;  (h]r�;  (hh e]r�;  (hhe]r�;  (hh	e]r�;  (h%heee]r�;  (ju*  ]r�;  (jw*  ]r�;  (jy*  ]r�;  (hh	e]r�;  (hh	e]r�;  (hjN  e]r�;  (j~*  ]r�;  (hhe]r�;  (hhe]r�;  (hjN  e]r�;  (j�-  ]r�;  (hh	e]r�;  (hh	eeee]r�;  (hh&ee]r�;  (h]r�;  (hh e]r�;  (hhe]r�;  (hh	e]r�;  (h%heeej�;  j�;  j�;  j�;  j�;  j�;  ]r�;  (ju*  ]r�;  (jw*  ]r�;  (jy*  ]r�;  (hh	e]r�;  (hh	e]r�;  (hjN  e]r�;  (j~*  ]r�;  (hh	e]r�;  (hhe]r�;  (hjN  e]r�;  (j�-  ]r�;  (hh	e]r�;  (hh	eeee]r�;  (hh&ee]r�;  (h]r�;  (hh e]r�;  (hhe]r�;  (hh	e]r�;  (h%heeej�;  j�;  j�;  j�;  ]r�;  (ju*  ]r�;  (jw*  ]r�;  (jy*  ]r�;  (hh	e]r�;  (hh	e]r�;  (hjN  e]r�;  (j~*  ]r�;  (hh	e]r�;  (hhe]r�;  (hjN  e]r�;  (j�-  ]r�;  (hh	e]r�;  (hh	eeee]r�;  (hh&ee]r�;  (h]r�;  (hh e]r�;  (hhe]r�;  (hh	e]r�;  (h%heeej�;  j�;  j�;  j�;  j�;  j�;  j�;  j�;  ]r�;  (ju*  ]r�;  (jw*  ]r�;  (jy*  ]r�;  (hh	e]r�;  (hh	e]r�;  (hjN  e]r�;  (j~*  ]r�;  (hh	e]r�;  (hhe]r�;  (hjN  e]r�;  (j�-  ]r�;  (hh	e]r�;  (hh	eeee]r�;  (hh&ee]r�;  (h]r�;  (hh e]r�;  (hhe]r�;  (hh	e]r�;  (h%heeej�;  j�;  ]r�;  (ju*  ]r�;  (jw*  ]r�;  (jy*  ]r�;  (hh	e]r�;  (hh	e]r�;  (hjN  e]r�;  (j~*  ]r�;  (hh	e]r�;  (hhe]r�;  (hjN  e]r�;  (j�-  ]r�;  (hh	e]r�;  (hh	eeee]r�;  (hh&ee]r�;  (h]r�;  (hh e]r�;  (hhe]r�;  (hh	e]r�;  (h%heeej�;  ]r�;  (ju*  ]r�;  (jw*  ]r�;  (jy*  ]r�;  (hh	e]r�;  (hh	e]r�;  (hjN  e]r�;  (j~*  ]r�;  (hh	e]r�;  (hhe]r�;  (hjN  e]r�;  (j�-  ]r�;  (hh	e]r�;  (hh	eeee]r�;  (hh&ee]r�;  (h]r�;  (hh e]r�;  (hhe]r�;  (hh	e]r�;  (h%heee]r�;  (ju*  ]r�;  (jw*  ]r <  (jy*  ]r<  (hh	e]r<  (hh	e]r<  (hjN  e]r<  (j~*  ]r<  (hh	e]r<  (hhe]r<  (hjN  e]r<  (j�-  ]r	<  (hh	e]r
<  (hh	eeee]r<  (hh&ee]r<  (h]r<  (hh e]r<  (hhe]r<  (hh	e]r<  (h%heee]r<  (ju*  ]r<  (jw*  ]r<  (jy*  ]r<  (hh	e]r<  (hh	e]r<  (hjN  e]r<  (j~*  ]r<  (hh	e]r<  (hhe]r<  (hjN  e]r<  (j�-  ]r<  (hh	e]r<  (hh	eeee]r<  (hh&ee]r<  (h]r <  (hh e]r!<  (hhe]r"<  (hh	e]r#<  (h%heeej<  ]r$<  (ju*  ]r%<  (jw*  ]r&<  (jy*  ]r'<  (hh	e]r(<  (hh	e]r)<  (hjN  e]r*<  (j~*  ]r+<  (hh	e]r,<  (hhe]r-<  (hjN  e]r.<  (j�-  ]r/<  (hh	e]r0<  (hh	eeee]r1<  (hh&ee]r2<  (h]r3<  (hh e]r4<  (hhe]r5<  (hh	e]r6<  (h%heeej$<  j$<  ]r7<  (ju*  ]r8<  (jw*  ]r9<  (jy*  ]r:<  (hh	e]r;<  (hh	e]r<<  (hjN  e]r=<  (j~*  ]r><  (hh	e]r?<  (hhe]r@<  (hjN  e]rA<  (j�-  ]rB<  (hh	e]rC<  (hh	eeee]rD<  (hh&ee]rE<  (h]rF<  (hh e]rG<  (hhe]rH<  (hhe]rI<  (h%heeej7<  ]rJ<  (ju*  ]rK<  (jw*  ]rL<  (jy*  ]rM<  (hh	e]rN<  (hh	e]rO<  (hjN  e]rP<  (j~*  ]rQ<  (hh	e]rR<  (hhe]rS<  (hjN  e]rT<  (j�-  ]rU<  (hh	e]rV<  (hh	eeee]rW<  (hh&ee]rX<  (h]rY<  (hh e]rZ<  (hhe]r[<  (hhe]r\<  (h%heeejJ<  ]r]<  (ju*  ]r^<  (jw*  ]r_<  (jy*  ]r`<  (hh	e]ra<  (hh	e]rb<  (hjN  e]rc<  (j~*  ]rd<  (hh	e]re<  (hhe]rf<  (hjN  e]rg<  (j�-  ]rh<  (hh	e]ri<  (hh	eeee]rj<  (hh&ee]rk<  (h]rl<  (hh e]rm<  (hhe]rn<  (hhe]ro<  (h%heeej]<  j]<  j]<  j]<  ]rp<  (ju*  ]rq<  (jw*  ]rr<  (jy*  ]rs<  (hh	e]rt<  (hh	e]ru<  (hjN  e]rv<  (j~*  ]rw<  (hh	e]rx<  (hhe]ry<  (hjN  e]rz<  (j�-  ]r{<  (hh	e]r|<  (hh	eeee]r}<  (hh&ee]r~<  (h]r<  (hh e]r�<  (hhe]r�<  (hhe]r�<  (h%heeejp<  ]r�<  (ju*  ]r�<  (jw*  ]r�<  (jy*  ]r�<  (hh	e]r�<  (hh	e]r�<  (hjN  e]r�<  (j~*  ]r�<  (hh	e]r�<  (hhe]r�<  (hjN  e]r�<  (j�-  ]r�<  (hh	e]r�<  (hh	eeee]r�<  (hh&ee]r�<  (h]r�<  (hh e]r�<  (hhe]r�<  (hhe]r�<  (h%heeej�<  j�<  j�<  ]r�<  (ju*  ]r�<  (jw*  ]r�<  (jy*  ]r�<  (hh	e]r�<  (hh	e]r�<  (hjN  e]r�<  (j~*  ]r�<  (hh	e]r�<  (hhe]r�<  (hjN  e]r�<  (j�-  ]r�<  (hh	e]r�<  (hh	eeee]r�<  (hh&ee]r�<  (h]r�<  (hh e]r�<  (hhe]r�<  (hhe]r�<  (h%heeej�<  j�<  j�<  j�<  j�<  ]r�<  (ju*  ]r�<  (jw*  ]r�<  (jy*  ]r�<  (hh	e]r�<  (hh	e]r�<  (hjN  e]r�<  (j~*  ]r�<  (hh	e]r�<  (hhe]r�<  (hjN  e]r�<  (j�-  ]r�<  (hh	e]r�<  (hh	eeee]r�<  (hh&ee]r�<  (h]r�<  (hh e]r�<  (hhe]r�<  (hhe]r�<  (h%heee]r�<  (ju*  ]r�<  (jw*  ]r�<  (jy*  ]r�<  (hh	e]r�<  (hh	e]r�<  (hjN  e]r�<  (j~*  ]r�<  (hhe]r�<  (hhe]r�<  (hjN  e]r�<  (j�-  ]r�<  (hh	e]r�<  (hh	eeee]r�<  (hh&ee]r�<  (h]r�<  (hh e]r�<  (hhe]r�<  (hhe]r�<  (h%heeej�<  ]r�<  (ju*  ]r�<  (jw*  ]r�<  (jy*  ]r�<  (hh	e]r�<  (hh	e]r�<  (hjN  e]r�<  (j~*  ]r�<  (hhe]r�<  (hhe]r�<  (hjN  e]r�<  (j�-  ]r�<  (hh	e]r�<  (hh	eeee]r�<  (hh&ee]r�<  (h]r�<  (hh e]r�<  (hhe]r�<  (hhe]r�<  (h%heeej�<  j�<  j�<  j�<  ]r�<  (ju*  ]r�<  (jw*  ]r�<  (jy*  ]r�<  (hh	e]r�<  (hh	e]r�<  (hjN  e]r�<  (j~*  ]r�<  (hhe]r�<  (hhe]r�<  (hjN  e]r�<  (j�-  ]r�<  (hh	e]r�<  (hh	eeee]r�<  (hh&ee]r�<  (h]r�<  (hh e]r�<  (hhe]r�<  (hhe]r�<  (h%heeej�<  j�<  j�<  j�<  ]r�<  (ju*  ]r�<  (jw*  ]r�<  (jy*  ]r�<  (hh	e]r�<  (hh	e]r�<  (hjN  e]r�<  (j~*  ]r�<  (hhe]r�<  (hhe]r�<  (hjN  e]r�<  (j�-  ]r =  (hh	e]r=  (hh	eeee]r=  (hh&ee]r=  (h]r=  (hh e]r=  (hhe]r=  (hhe]r=  (h%heeej�<  j�<  j�<  j�<  j�<  ]r=  (ju*  ]r	=  (jw*  ]r
=  (jy*  ]r=  (hh	e]r=  (hh	e]r=  (hjN  e]r=  (j~*  ]r=  (hhe]r=  (hhe]r=  (hjN  e]r=  (j�-  ]r=  (hh	e]r=  (hh	eeee]r=  (hh&ee]r=  (h]r=  (hh e]r=  (hhe]r=  (hhe]r=  (h%heeej=  ]r=  (ju*  ]r=  (jw*  ]r=  (jy*  ]r=  (hh	e]r=  (hh	e]r =  (hjN  e]r!=  (j~*  ]r"=  (hhe]r#=  (hhe]r$=  (hjN  e]r%=  (j�-  ]r&=  (hh	e]r'=  (hh	eeee]r(=  (hh&ee]r)=  (h]r*=  (hh e]r+=  (hhe]r,=  (hhe]r-=  (h%heeej=  j=  j=  j=  j=  j=  j=  j=  j=  ]r.=  (ju*  ]r/=  (jw*  ]r0=  (jy*  ]r1=  (hh	e]r2=  (hh	e]r3=  (hjN  e]r4=  (j~*  ]r5=  (hhe]r6=  (hhe]r7=  (hjN  e]r8=  (j�-  ]r9=  (hh	e]r:=  (hh	eeee]r;=  (hh&ee]r<=  (h]r==  (hh e]r>=  (hhe]r?=  (hhe]r@=  (h%heeej.=  j.=  j.=  j.=  j.=  j.=  j.=  ]rA=  (ju*  ]rB=  (jw*  ]rC=  (jy*  ]rD=  (hh	e]rE=  (hh	e]rF=  (hjN  e]rG=  (j~*  ]rH=  (hhe]rI=  (hhe]rJ=  (hjN  e]rK=  (j�-  ]rL=  (hh	e]rM=  (hh	eeee]rN=  (hh&ee]rO=  (h]rP=  (hh e]rQ=  (hhe]rR=  (hhe]rS=  (h%heeejA=  ]rT=  (ju*  ]rU=  (jw*  ]rV=  (jy*  ]rW=  (hh	e]rX=  (hh	e]rY=  (hjN  e]rZ=  (j~*  ]r[=  (hhe]r\=  (hhe]r]=  (hjN  e]r^=  (j�-  ]r_=  (hh	e]r`=  (hh	eeee]ra=  (hh&ee]rb=  (h]rc=  (hh e]rd=  (hhe]re=  (hhe]rf=  (h%heeejT=  jT=  ]rg=  (ju*  ]rh=  (jw*  ]ri=  (jy*  ]rj=  (hh	e]rk=  (hh	e]rl=  (hjN  e]rm=  (j~*  ]rn=  (hhe]ro=  (hhe]rp=  (hjN  e]rq=  (j�-  ]rr=  (hh	e]rs=  (hh	eeee]rt=  (hh&ee]ru=  (h]rv=  (hh e]rw=  (hhe]rx=  (hhe]ry=  (h%heee]rz=  (ju*  ]r{=  (jw*  ]r|=  (jy*  ]r}=  (hh	e]r~=  (hh	e]r=  (hjN  e]r�=  (j~*  ]r�=  (hhe]r�=  (hhe]r�=  (hjN  e]r�=  (j�-  ]r�=  (hh	e]r�=  (hh	eeee]r�=  (hh&ee]r�=  (h]r�=  (hh e]r�=  (hhe]r�=  (hhe]r�=  (h%heee]r�=  (ju*  ]r�=  (jw*  ]r�=  (jy*  ]r�=  (hh	e]r�=  (hh	e]r�=  (hjN  e]r�=  (j~*  ]r�=  (hhe]r�=  (hhe]r�=  (hjN  e]r�=  (j�-  ]r�=  (hh	e]r�=  (hh	eeee]r�=  (hh&ee]r�=  (h]r�=  (hh e]r�=  (hhe]r�=  (hhe]r�=  (h%heeej�=  e(]r�=  (X   Normsr�=  ]r�=  (X   Oblr�=  ]r�=  (X   Movedr�=  ]r�=  (hh	e]r�=  (hj�)  e]r�=  (hjN  e]r�=  (X   Movedr�=  ]r�=  (hh	e]r�=  (hj�)  e]r�=  (hh&e]r�=  (X	   Next-Mover�=  ]r�=  (hh	e]r�=  (hh	eeee]r�=  (hhee]r�=  (h]r�=  (hh e]r�=  (hh	e]r�=  (hhe]r�=  (h%h&eeej�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  ]r�=  (j�=  ]r�=  (j�=  ]r�=  (j�=  ]r�=  (hh	e]r�=  (hj�)  e]r�=  (hjN  e]r�=  (j�=  ]r�=  (hh	e]r�=  (hj�)  e]r�=  (hh&e]r�=  (j�=  ]r�=  (hh	e]r�=  (hh	eeee]r�=  (hhee]r�=  (h]r�=  (hh e]r�=  (hh	e]r�=  (hhe]r�=  (h%h&eeej�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  ]r�=  (j�=  ]r�=  (j�=  ]r�=  (j�=  ]r�=  (hh	e]r�=  (hj�)  e]r�=  (hjN  e]r�=  (j�=  ]r�=  (hh	e]r�=  (hj�)  e]r�=  (hh&e]r�=  (j�=  ]r�=  (hh	e]r�=  (hh	eeee]r�=  (hhee]r�=  (h]r�=  (hh e]r�=  (hh	e]r�=  (hhe]r�=  (h%h&eeej�=  j�=  j�=  j�=  ]r�=  (j�=  ]r�=  (j�=  ]r�=  (j�=  ]r�=  (hh	e]r�=  (hj�)  e]r�=  (hjN  e]r�=  (j�=  ]r�=  (hh	e]r�=  (hj�)  e]r�=  (hh&e]r�=  (j�=  ]r�=  (hh	e]r�=  (hh	eeee]r�=  (hhee]r�=  (h]r�=  (hh e]r�=  (hh	e]r�=  (hhe]r�=  (h%h&eeej�=  ]r�=  (j�=  ]r�=  (j�=  ]r�=  (j�=  ]r�=  (hh	e]r�=  (hj�)  e]r�=  (hjN  e]r�=  (j�=  ]r�=  (hh	e]r�=  (hj�)  e]r�=  (hh&e]r�=  (j�=  ]r�=  (hh	e]r�=  (hh	eeee]r�=  (hhee]r�=  (h]r >  (hh e]r>  (hh	e]r>  (hhe]r>  (h%h&eee]r>  (j�=  ]r>  (j�=  ]r>  (j�=  ]r>  (hh	e]r>  (hj�)  e]r	>  (hjN  e]r
>  (j�=  ]r>  (hh	e]r>  (hj�)  e]r>  (hh&e]r>  (j�=  ]r>  (hh	e]r>  (hh	eeee]r>  (hhee]r>  (h]r>  (hh e]r>  (hh	e]r>  (hhe]r>  (h%h&eeej>  j>  j>  j>  j>  j>  ]r>  (j�=  ]r>  (j�=  ]r>  (j�=  ]r>  (hh	e]r>  (hj�)  e]r>  (hjN  e]r>  (j�=  ]r>  (hh	e]r>  (hj�)  e]r >  (hh&e]r!>  (j�=  ]r">  (hh	e]r#>  (hh	eeee]r$>  (hhee]r%>  (h]r&>  (hh e]r'>  (hh	e]r(>  (hhe]r)>  (h%h&eeej>  j>  ]r*>  (j�=  ]r+>  (j�=  ]r,>  (j�=  ]r->  (hh	e]r.>  (hj�)  e]r/>  (hjN  e]r0>  (j�=  ]r1>  (hh	e]r2>  (hj�)  e]r3>  (hh&e]r4>  (j�=  ]r5>  (hh	e]r6>  (hh	eeee]r7>  (hhee]r8>  (h]r9>  (hh e]r:>  (hh	e]r;>  (hhe]r<>  (h%h&eeej*>  j*>  j*>  j*>  j*>  j*>  j*>  j*>  j*>  ]r=>  (j�=  ]r>>  (j�=  ]r?>  (j�=  ]r@>  (hh	e]rA>  (hj�)  e]rB>  (hjN  e]rC>  (j�=  ]rD>  (hh	e]rE>  (hj�)  e]rF>  (hh&e]rG>  (j�=  ]rH>  (hh	e]rI>  (hh	eeee]rJ>  (hhee]rK>  (h]rL>  (hh e]rM>  (hh	e]rN>  (hhe]rO>  (h%h&eeej=>  ]rP>  (j�=  ]rQ>  (j�=  ]rR>  (j�=  ]rS>  (hh	e]rT>  (hj�)  e]rU>  (hjN  e]rV>  (j�=  ]rW>  (hh	e]rX>  (hj�)  e]rY>  (hh&e]rZ>  (j�=  ]r[>  (hh	e]r\>  (hh	eeee]r]>  (hhee]r^>  (h]r_>  (hh e]r`>  (hh	e]ra>  (hhe]rb>  (h%h&eeejP>  jP>  ]rc>  (j�=  ]rd>  (j�=  ]re>  (j�=  ]rf>  (hh	e]rg>  (hj�)  e]rh>  (hjN  e]ri>  (j�=  ]rj>  (hh	e]rk>  (hj�)  e]rl>  (hh&e]rm>  (j�=  ]rn>  (hh	e]ro>  (hh	eeee]rp>  (hhee]rq>  (h]rr>  (hh e]rs>  (hh	e]rt>  (hhe]ru>  (h%h&eee]rv>  (j�=  ]rw>  (j�=  ]rx>  (j�=  ]ry>  (hh	e]rz>  (hj�)  e]r{>  (hjN  e]r|>  (j�=  ]r}>  (hh	e]r~>  (hj�)  e]r>  (hh&e]r�>  (j�=  ]r�>  (hh	e]r�>  (hh	eeee]r�>  (hhee]r�>  (h]r�>  (hh e]r�>  (hh	e]r�>  (hhe]r�>  (h%h&eeejv>  jv>  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (hh	e]r�>  (hj�)  e]r�>  (hjN  e]r�>  (j�=  ]r�>  (hh	e]r�>  (hj�)  e]r�>  (hh&e]r�>  (j�=  ]r�>  (hh	e]r�>  (hh	eeee]r�>  (hhee]r�>  (h]r�>  (hh e]r�>  (hh	e]r�>  (hhe]r�>  (h%h&eeej�>  j�>  j�>  j�>  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (hh	e]r�>  (hj�)  e]r�>  (hjN  e]r�>  (j�=  ]r�>  (hh	e]r�>  (hj�)  e]r�>  (hh&e]r�>  (j�=  ]r�>  (hh	e]r�>  (hh	eeee]r�>  (hhee]r�>  (h]r�>  (hh e]r�>  (hh	e]r�>  (hhe]r�>  (h%h&eeej�>  j�>  j�>  j�>  j�>  j�>  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (hh	e]r�>  (hj�)  e]r�>  (hjN  e]r�>  (j�=  ]r�>  (hh	e]r�>  (hj�)  e]r�>  (hh&e]r�>  (j�=  ]r�>  (hh	e]r�>  (hh	eeee]r�>  (hhee]r�>  (h]r�>  (hh e]r�>  (hh	e]r�>  (hhe]r�>  (h%h&eeej�>  j�>  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (hh	e]r�>  (hj�)  e]r�>  (hjN  e]r�>  (j�=  ]r�>  (hh	e]r�>  (hj�)  e]r�>  (hh&e]r�>  (j�=  ]r�>  (hh	e]r�>  (hh	eeee]r�>  (hhee]r�>  (h]r�>  (hh e]r�>  (hh	e]r�>  (hhe]r�>  (h%h&eee]r�>  (j�=  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (hh	e]r�>  (hj�)  e]r�>  (hjN  e]r�>  (j�=  ]r�>  (hh	e]r�>  (hj�)  e]r�>  (hh&e]r�>  (j�=  ]r�>  (hh	e]r�>  (hh	eeee]r�>  (hhee]r�>  (h]r�>  (hh e]r�>  (hh	e]r�>  (hhe]r�>  (h%h&eeej�>  j�>  j�>  j�>  j�>  j�>  j�>  j�>  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (hj�)  e]r�>  (hj�)  e]r�>  (hjN  e]r�>  (j�=  ]r�>  (hh	e]r�>  (hj�)  e]r�>  (hh&e]r�>  (j�=  ]r�>  (hh	e]r�>  (hh	eeee]r�>  (hhee]r�>  (h]r�>  (hh e]r�>  (hh	e]r�>  (hhe]r�>  (h%h&eeej�>  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (j�=  ]r�>  (hj�)  e]r�>  (hj�)  e]r ?  (hjN  e]r?  (j�=  ]r?  (hh	e]r?  (hj�)  e]r?  (hh&e]r?  (j�=  ]r?  (hh	e]r?  (hh	eeee]r?  (hhee]r	?  (h]r
?  (hh e]r?  (hh	e]r?  (hhe]r?  (h%h&eeej�>  j�>  j�>  ]r?  (j�=  ]r?  (j�=  ]r?  (j�=  ]r?  (hh	e]r?  (hj�)  e]r?  (hjN  e]r?  (j�=  ]r?  (hh	e]r?  (hj�)  e]r?  (hh&e]r?  (j�=  ]r?  (hh	e]r?  (hh	eeee]r?  (hhee]r?  (h]r?  (hh e]r?  (hh	e]r?  (hhe]r ?  (h%h&eee]r!?  (j�=  ]r"?  (j�=  ]r#?  (j�=  ]r$?  (hh	e]r%?  (hj�)  e]r&?  (hjN  e]r'?  (j�=  ]r(?  (hh	e]r)?  (hj�)  e]r*?  (hh&e]r+?  (j�=  ]r,?  (hh	e]r-?  (hh	eeee]r.?  (hhee]r/?  (h]r0?  (hh e]r1?  (hh	e]r2?  (hhe]r3?  (h%h&eee]r4?  (j�=  ]r5?  (j�=  ]r6?  (j�=  ]r7?  (hh	e]r8?  (hj�)  e]r9?  (hjN  e]r:?  (j�=  ]r;?  (hh	e]r<?  (hj�)  e]r=?  (hh&e]r>?  (j�=  ]r??  (hh	e]r@?  (hh	eeee]rA?  (hhee]rB?  (h]rC?  (hh e]rD?  (hh	e]rE?  (hhe]rF?  (h%h&eeej4?  j4?  j4?  j4?  j4?  j4?  j4?  j4?  ]rG?  (j�=  ]rH?  (j�=  ]rI?  (j�=  ]rJ?  (hh	e]rK?  (hj�)  e]rL?  (hjN  e]rM?  (j�=  ]rN?  (hh	e]rO?  (hj�)  e]rP?  (hh&e]rQ?  (j�=  ]rR?  (hh	e]rS?  (hh	eeee]rT?  (hhee]rU?  (h]rV?  (hh e]rW?  (hh	e]rX?  (hhe]rY?  (h%h&eeejG?  jG?  ]rZ?  (j�=  ]r[?  (j�=  ]r\?  (j�=  ]r]?  (hh	e]r^?  (hj�)  e]r_?  (hjN  e]r`?  (j�=  ]ra?  (hj�)  e]rb?  (hj�)  e]rc?  (hh&e]rd?  (j�=  ]re?  (hh	e]rf?  (hh	eeee]rg?  (hhee]rh?  (h]ri?  (hh e]rj?  (hh	e]rk?  (hhe]rl?  (h%h&eeejZ?  jZ?  jZ?  jZ?  ]rm?  (j�=  ]rn?  (j�=  ]ro?  (j�=  ]rp?  (hh	e]rq?  (hj�)  e]rr?  (hjN  e]rs?  (j�=  ]rt?  (hj�)  e]ru?  (hj�)  e]rv?  (hh&e]rw?  (j�=  ]rx?  (hh	e]ry?  (hh	eeee]rz?  (hhee]r{?  (h]r|?  (hh e]r}?  (hh	e]r~?  (hhe]r?  (h%h&eee]r�?  (j�=  ]r�?  (j�=  ]r�?  (j�=  ]r�?  (hh	e]r�?  (hj�)  e]r�?  (hjN  e]r�?  (j�=  ]r�?  (hj�)  e]r�?  (hj�)  e]r�?  (hh&e]r�?  (X	   Next-Mover�?  ]r�?  (hh	e]r�?  (hh	eeee]r�?  (hhee]r�?  (h]r�?  (hh e]r�?  (hh	e]r�?  (hhe]r�?  (h%h&eee]r�?  (j�=  ]r�?  (j�=  ]r�?  (j�=  ]r�?  (hh	e]r�?  (hj�)  e]r�?  (hjN  e]r�?  (j�=  ]r�?  (hj�)  e]r�?  (hj�)  e]r�?  (hh&e]r�?  (j�?  ]r�?  (hh	e]r�?  (hh	eeee]r�?  (hhee]r�?  (h]r�?  (hh e]r�?  (hh	e]r�?  (hhe]r�?  (h%h&eee]r�?  (j�=  ]r�?  (j�=  ]r�?  (j�=  ]r�?  (hh	e]r�?  (hj�)  e]r�?  (hjN  e]r�?  (j�=  ]r�?  (hj�)  e]r�?  (hj�)  e]r�?  (hh&e]r�?  (j�?  ]r�?  (hh	e]r�?  (hh	eeee]r�?  (hhee]r�?  (h]r�?  (hh e]r�?  (hh	e]r�?  (hhe]r�?  (h%h&eeej�?  ]r�?  (j�=  ]r�?  (j�=  ]r�?  (j�=  ]r�?  (hh	e]r�?  (hj�)  e]r�?  (hjN  e]r�?  (j�=  ]r�?  (hj�)  e]r�?  (hj�)  e]r�?  (hh&e]r�?  (j�?  ]r�?  (hh	e]r�?  (hh	eeee]r�?  (hhee]r�?  (h]r�?  (hh e]r�?  (hh	e]r�?  (hhe]r�?  (h%h&eeej�?  ]r�?  (j�=  ]r�?  (j�=  ]r�?  (j�=  ]r�?  (hh	e]r�?  (hj�)  e]r�?  (hjN  e]r�?  (j�=  ]r�?  (hj�)  e]r�?  (hj�)  e]r�?  (hh&e]r�?  (j�?  ]r�?  (hh	e]r�?  (hh	eeee]r�?  (hhee]r�?  (h]r�?  (hh e]r�?  (hh	e]r�?  (hhe]r�?  (h%h&eee]r�?  (j�=  ]r�?  (j�=  ]r�?  (j�=  ]r�?  (hh	e]r�?  (hj�)  e]r�?  (hjN  e]r�?  (j�=  ]r�?  (hj�)  e]r�?  (hj�)  e]r�?  (hh&e]r�?  (j�?  ]r�?  (hh	e]r�?  (hh	eeee]r�?  (hhee]r�?  (h]r�?  (hh e]r�?  (hh	e]r�?  (hhe]r�?  (h%h&eeej�?  j�?  j�?  j�?  j�?  j�?  j�?  j�?  j�?  ]r�?  (j�=  ]r�?  (j�=  ]r�?  (j�=  ]r�?  (hh	e]r�?  (hj�)  e]r�?  (hjN  e]r�?  (j�=  ]r�?  (hj�)  e]r�?  (hj�)  e]r�?  (hh&e]r�?  (j�?  ]r�?  (hh	e]r�?  (hh	eeee]r @  (hhee]r@  (h]r@  (hh e]r@  (hh	e]r@  (hhe]r@  (h%h&eeej�?  ]r@  (j�=  ]r@  (j�=  ]r@  (j�=  ]r	@  (hh	e]r
@  (hj�)  e]r@  (hjN  e]r@  (j�=  ]r@  (hj�)  e]r@  (hj�)  e]r@  (hh&e]r@  (j�?  ]r@  (hh	e]r@  (hh	eeee]r@  (hhee]r@  (h]r@  (hh e]r@  (hh	e]r@  (hhe]r@  (h%h&eeej@  j@  j@  j@  ]r@  (j�=  ]r@  (j�=  ]r@  (j�=  ]r@  (hh	e]r@  (hj�)  e]r@  (hjN  e]r@  (j�=  ]r @  (hj�)  e]r!@  (hj�)  e]r"@  (hh&e]r#@  (j�?  ]r$@  (hh	e]r%@  (hh	eeee]r&@  (hhee]r'@  (h]r(@  (hh e]r)@  (hh	e]r*@  (hhe]r+@  (h%h&eeej@  j@  j@  j@  j@  ]r,@  (j�=  ]r-@  (j�=  ]r.@  (j�=  ]r/@  (hh	e]r0@  (hj�)  e]r1@  (hjN  e]r2@  (j�=  ]r3@  (hj�)  e]r4@  (hj�)  e]r5@  (hh&e]r6@  (j�?  ]r7@  (hh	e]r8@  (hh	eeee]r9@  (hhee]r:@  (h]r;@  (hh e]r<@  (hh	e]r=@  (hhe]r>@  (h%h&eeej,@  j,@  j,@  j,@  j,@  j,@  j,@  j,@  j,@  ]r?@  (j�=  ]r@@  (j�=  ]rA@  (j�=  ]rB@  (hh	e]rC@  (hj�)  e]rD@  (hjN  e]rE@  (j�=  ]rF@  (hh	e]rG@  (hj�)  e]rH@  (hh&e]rI@  (j�?  ]rJ@  (hh	e]rK@  (hh	eeee]rL@  (hhee]rM@  (h]rN@  (hh e]rO@  (hh	e]rP@  (hhe]rQ@  (h%h&eeej?@  j?@  ]rR@  (j�=  ]rS@  (j�=  ]rT@  (j�=  ]rU@  (hh	e]rV@  (hj�)  e]rW@  (hjN  e]rX@  (j�=  ]rY@  (hh	e]rZ@  (hj�)  e]r[@  (hh&e]r\@  (j�?  ]r]@  (hh	e]r^@  (hh	eeee]r_@  (hhee]r`@  (h]ra@  (hh e]rb@  (hh	e]rc@  (hhe]rd@  (h%h&eee]re@  (j�=  ]rf@  (j�=  ]rg@  (j�=  ]rh@  (hh	e]ri@  (hj�)  e]rj@  (hjN  e]rk@  (j�=  ]rl@  (hh	e]rm@  (hj�)  e]rn@  (hh&e]ro@  (j�?  ]rp@  (hh	e]rq@  (hh	eeee]rr@  (hhee]rs@  (h]rt@  (hh e]ru@  (hh	e]rv@  (hhe]rw@  (h%h&eee]rx@  (j�=  ]ry@  (j�=  ]rz@  (j�=  ]r{@  (hh	e]r|@  (hj�)  e]r}@  (hjN  e]r~@  (j�=  ]r@  (hh	e]r�@  (hj�)  e]r�@  (hh&e]r�@  (j�?  ]r�@  (hh	e]r�@  (hh	eeee]r�@  (hhee]r�@  (h]r�@  (hh e]r�@  (hh	e]r�@  (hhe]r�@  (h%h&eeejx@  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (hh	e]r�@  (hj�)  e]r�@  (hjN  e]r�@  (j�=  ]r�@  (hh	e]r�@  (hj�)  e]r�@  (hh&e]r�@  (j�?  ]r�@  (hh	e]r�@  (hh	eeee]r�@  (hhee]r�@  (h]r�@  (hh e]r�@  (hh	e]r�@  (hhe]r�@  (h%h&eeej�@  j�@  j�@  j�@  j�@  j�@  j�@  j�@  j�@  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (hh	e]r�@  (hj�)  e]r�@  (hjN  e]r�@  (j�=  ]r�@  (hj�)  e]r�@  (hj�)  e]r�@  (hh&e]r�@  (j�?  ]r�@  (hh	e]r�@  (hh	eeee]r�@  (hhee]r�@  (h]r�@  (hh e]r�@  (hh	e]r�@  (hhe]r�@  (h%h&eeej�@  j�@  j�@  j�@  j�@  j�@  j�@  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (hh	e]r�@  (hj�)  e]r�@  (hjN  e]r�@  (j�=  ]r�@  (hj�)  e]r�@  (hj�)  e]r�@  (hh&e]r�@  (j�?  ]r�@  (hh	e]r�@  (hh	eeee]r�@  (hhee]r�@  (h]r�@  (hh e]r�@  (hh	e]r�@  (hhe]r�@  (h%h&eeej�@  j�@  j�@  j�@  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (hh	e]r�@  (hj�)  e]r�@  (hjN  e]r�@  (j�=  ]r�@  (hj�)  e]r�@  (hj�)  e]r�@  (hh&e]r�@  (j�?  ]r�@  (hh	e]r�@  (hh	eeee]r�@  (hhee]r�@  (h]r�@  (hh e]r�@  (hh	e]r�@  (hhe]r�@  (h%h&eeej�@  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (hj�)  e]r�@  (hj�)  e]r�@  (hjN  e]r�@  (j�=  ]r�@  (hj�)  e]r�@  (hj�)  e]r�@  (hh&e]r�@  (j�?  ]r�@  (hh	e]r�@  (hh	eeee]r�@  (hhee]r�@  (h]r�@  (hh e]r�@  (hh	e]r�@  (hhe]r�@  (h%h&eeej�@  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (hj�)  e]r�@  (hj�)  e]r�@  (hjN  e]r�@  (j�=  ]r�@  (hj�)  e]r�@  (hj�)  e]r�@  (hh&e]r�@  (j�?  ]r�@  (hh	e]r�@  (hh	eeee]r�@  (hhee]r�@  (h]r�@  (hh e]r�@  (hh	e]r�@  (hhe]r�@  (h%h&eeej�@  j�@  ]r�@  (j�=  ]r�@  (j�=  ]r�@  (j�=  ]r A  (hj�)  e]rA  (hj�)  e]rA  (hjN  e]rA  (j�=  ]rA  (hj�)  e]rA  (hj�)  e]rA  (hh&e]rA  (j�?  ]rA  (hh	e]r	A  (hh	eeee]r
A  (hhee]rA  (h]rA  (hh e]rA  (hh	e]rA  (hhe]rA  (h%h&eeej�@  j�@  ]rA  (j�=  ]rA  (j�=  ]rA  (j�=  ]rA  (hj�)  e]rA  (hj�)  e]rA  (hjN  e]rA  (j�=  ]rA  (hj�)  e]rA  (hj�)  e]rA  (hh&e]rA  (j�?  ]rA  (hh	e]rA  (hh	eeee]rA  (hhee]rA  (h]rA  (hh e]r A  (hh	e]r!A  (hhe]r"A  (h%h&eee]r#A  (j�=  ]r$A  (j�=  ]r%A  (j�=  ]r&A  (hj�)  e]r'A  (hj�)  e]r(A  (hjN  e]r)A  (j�=  ]r*A  (hh	e]r+A  (hj�)  e]r,A  (hh&e]r-A  (j�?  ]r.A  (hh	e]r/A  (hh	eeee]r0A  (hhee]r1A  (h]r2A  (hh e]r3A  (hh	e]r4A  (hhe]r5A  (h%h&eee]r6A  (j�=  ]r7A  (j�=  ]r8A  (j�=  ]r9A  (hj�)  e]r:A  (hj�)  e]r;A  (hjN  e]r<A  (j�=  ]r=A  (hh	e]r>A  (hj�)  e]r?A  (hh&e]r@A  (j�?  ]rAA  (hh	e]rBA  (hh	eeee]rCA  (hhee]rDA  (h]rEA  (hh e]rFA  (hh	e]rGA  (hhe]rHA  (h%h&eeej6A  j6A  j6A  j6A  j6A  j6A  ]rIA  (j�=  ]rJA  (j�=  ]rKA  (j�=  ]rLA  (hj�)  e]rMA  (hj�)  e]rNA  (hjN  e]rOA  (j�=  ]rPA  (hh	e]rQA  (hj�)  e]rRA  (hh&e]rSA  (j�?  ]rTA  (hh	e]rUA  (hh	eeee]rVA  (hhee]rWA  (h]rXA  (hh e]rYA  (hh	e]rZA  (hhe]r[A  (h%h&eeejIA  jIA  ]r\A  (j�=  ]r]A  (j�=  ]r^A  (j�=  ]r_A  (hj�)  e]r`A  (hj�)  e]raA  (hjN  e]rbA  (j�=  ]rcA  (hh	e]rdA  (hj�)  e]reA  (hh&e]rfA  (j�?  ]rgA  (hh	e]rhA  (hh	eeee]riA  (hhee]rjA  (h]rkA  (hh e]rlA  (hh	e]rmA  (hhe]rnA  (h%h&eee]roA  (j�=  ]rpA  (j�=  ]rqA  (j�=  ]rrA  (hj�)  e]rsA  (hj�)  e]rtA  (hjN  e]ruA  (j�=  ]rvA  (hh	e]rwA  (hj�)  e]rxA  (hh&e]ryA  (j�?  ]rzA  (hh	e]r{A  (hh	eeee]r|A  (hhee]r}A  (h]r~A  (hh e]rA  (hh	e]r�A  (hhe]r�A  (h%h&eee]r�A  (j�=  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (hj�)  e]r�A  (hj�)  e]r�A  (hjN  e]r�A  (j�=  ]r�A  (hh	e]r�A  (hj�)  e]r�A  (hh&e]r�A  (j�?  ]r�A  (hh	e]r�A  (hh	eeee]r�A  (hhee]r�A  (h]r�A  (hh e]r�A  (hh	e]r�A  (hhe]r�A  (h%h&eeej�A  j�A  j�A  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (hj�)  e]r�A  (hj�)  e]r�A  (hjN  e]r�A  (j�=  ]r�A  (hh	e]r�A  (hj�)  e]r�A  (hh&e]r�A  (j�?  ]r�A  (hh	e]r�A  (hh	eeee]r�A  (hhee]r�A  (h]r�A  (hh e]r�A  (hh	e]r�A  (hhe]r�A  (h%h&eeej�A  j�A  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (hj�)  e]r�A  (hj�)  e]r�A  (hjN  e]r�A  (j�=  ]r�A  (hh	e]r�A  (hj�)  e]r�A  (hh&e]r�A  (j�?  ]r�A  (hh	e]r�A  (hh	eeee]r�A  (hhee]r�A  (h]r�A  (hh e]r�A  (hh	e]r�A  (hhe]r�A  (h%h&eeej�A  j�A  j�A  j�A  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (hj�)  e]r�A  (hj�)  e]r�A  (hjN  e]r�A  (j�=  ]r�A  (hh	e]r�A  (hj�)  e]r�A  (hh&e]r�A  (j�?  ]r�A  (hh	e]r�A  (hh	eeee]r�A  (hhee]r�A  (h]r�A  (hh e]r�A  (hh	e]r�A  (hhe]r�A  (h%h&eee]r�A  (j�=  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (hj�)  e]r�A  (hj�)  e]r�A  (hjN  e]r�A  (j�=  ]r�A  (hh	e]r�A  (hj�)  e]r�A  (hh&e]r�A  (j�?  ]r�A  (hh	e]r�A  (hh	eeee]r�A  (hhee]r�A  (h]r�A  (hh e]r�A  (hh	e]r�A  (hhe]r�A  (h%h&eeej�A  j�A  j�A  j�A  j�A  j�A  j�A  j�A  j�A  j�A  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (hj�)  e]r�A  (hj�)  e]r�A  (hjN  e]r�A  (j�=  ]r�A  (hh	e]r�A  (hj�)  e]r�A  (hh&e]r�A  (j�?  ]r�A  (hh	e]r�A  (hh	eeee]r�A  (hhee]r�A  (h]r�A  (hh e]r�A  (hh	e]r�A  (hhe]r�A  (h%h&eeej�A  j�A  j�A  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (j�=  ]r�A  (hj�)  e]r�A  (hj�)  e]r�A  (hjN  e]r�A  (j�=  ]r�A  (hh	e]r�A  (hj�)  e]r�A  (hh&e]r�A  (j�?  ]r�A  (hh	e]r B  (hh	eeee]rB  (hhee]rB  (h]rB  (hh e]rB  (hh	e]rB  (hhe]rB  (h%h&eee]rB  (j�=  ]rB  (j�=  ]r	B  (j�=  ]r
B  (hj�)  e]rB  (hj�)  e]rB  (hjN  e]rB  (j�=  ]rB  (hh	e]rB  (hj�)  e]rB  (hh&e]rB  (j�?  ]rB  (hh	e]rB  (hh	eeee]rB  (hhee]rB  (h]rB  (hh e]rB  (hh	e]rB  (hhe]rB  (h%h&eeejB  jB  ]rB  (j�=  ]rB  (j�=  ]rB  (j�=  ]rB  (hj�)  e]rB  (hj�)  e]rB  (hjN  e]r B  (j�=  ]r!B  (hh	e]r"B  (hj�)  e]r#B  (hh&e]r$B  (j�?  ]r%B  (hh	e]r&B  (hh	eeee]r'B  (hhee]r(B  (h]r)B  (hh e]r*B  (hh	e]r+B  (hhe]r,B  (h%h&eeejB  jB  jB  ]r-B  (j�=  ]r.B  (j�=  ]r/B  (j�=  ]r0B  (hj�)  e]r1B  (hj�)  e]r2B  (hjN  e]r3B  (j�=  ]r4B  (hh	e]r5B  (hj�)  e]r6B  (hh&e]r7B  (j�?  ]r8B  (hh	e]r9B  (hh	eeee]r:B  (hhee]r;B  (h]r<B  (hh e]r=B  (hh	e]r>B  (hhe]r?B  (h%h&eeej-B  j-B  j-B  j-B  j-B  ]r@B  (j�=  ]rAB  (j�=  ]rBB  (j�=  ]rCB  (hh	e]rDB  (hj�)  e]rEB  (hjN  e]rFB  (j�=  ]rGB  (hh	e]rHB  (hj�)  e]rIB  (hh&e]rJB  (j�?  ]rKB  (hh	e]rLB  (hh	eeee]rMB  (hhee]rNB  (h]rOB  (hh e]rPB  (hh	e]rQB  (hhe]rRB  (h%h&eeej@B  ]rSB  (j�=  ]rTB  (j�=  ]rUB  (j�=  ]rVB  (hh	e]rWB  (hj�)  e]rXB  (hjN  e]rYB  (j�=  ]rZB  (hh	e]r[B  (hj�)  e]r\B  (hh&e]r]B  (j�?  ]r^B  (hh	e]r_B  (hh	eeee]r`B  (hhee]raB  (h]rbB  (hh e]rcB  (hh	e]rdB  (hhe]reB  (h%h&eeejSB  jSB  jSB  jSB  jSB  jSB  jSB  jSB  ]rfB  (j�=  ]rgB  (j�=  ]rhB  (j�=  ]riB  (hh	e]rjB  (hj�)  e]rkB  (hjN  e]rlB  (j�=  ]rmB  (hh	e]rnB  (hj�)  e]roB  (hh&e]rpB  (j�?  ]rqB  (hh	e]rrB  (hh	eeee]rsB  (hhee]rtB  (h]ruB  (hh e]rvB  (hh	e]rwB  (hhe]rxB  (h%h&eee]ryB  (j�=  ]rzB  (j�=  ]r{B  (j�=  ]r|B  (hh	e]r}B  (hj�)  e]r~B  (hjN  e]rB  (j�=  ]r�B  (hh	e]r�B  (hj�)  e]r�B  (hh&e]r�B  (j�?  ]r�B  (hh	e]r�B  (hh	eeee]r�B  (hhee]r�B  (h]r�B  (hh e]r�B  (hh	e]r�B  (hhe]r�B  (h%h&eeejyB  ]r�B  (j�=  ]r�B  (j�=  ]r�B  (j�=  ]r�B  (hj�)  e]r�B  (hj�)  e]r�B  (hjN  e]r�B  (j�=  ]r�B  (hh	e]r�B  (hj�)  e]r�B  (hh&e]r�B  (j�?  ]r�B  (hh	e]r�B  (hh	eeee]r�B  (hhee]r�B  (h]r�B  (hh e]r�B  (hh	e]r�B  (hhe]r�B  (h%h&eeej�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  ]r�B  (j�=  ]r�B  (j�=  ]r�B  (j�=  ]r�B  (hj�)  e]r�B  (hj�)  e]r�B  (hjN  e]r�B  (j�=  ]r�B  (hh	e]r�B  (hj�)  e]r�B  (hh&e]r�B  (j�?  ]r�B  (hh	e]r�B  (hh	eeee]r�B  (hhee]r�B  (h]r�B  (hh e]r�B  (hh	e]r�B  (hhe]r�B  (h%h&eeej�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  ]r�B  (j�=  ]r�B  (j�=  ]r�B  (j�=  ]r�B  (hj�)  e]r�B  (hj�)  e]r�B  (hjN  e]r�B  (j�=  ]r�B  (hh	e]r�B  (hj�)  e]r�B  (hh&e]r�B  (j�?  ]r�B  (hh	e]r�B  (hh	eeee]r�B  (hhee]r�B  (h]r�B  (hh e]r�B  (hh	e]r�B  (hhe]r�B  (h%h&eeej�B  ]r�B  (j�=  ]r�B  (j�=  ]r�B  (j�=  ]r�B  (hj�)  e]r�B  (hj�)  e]r�B  (hjN  e]r�B  (j�=  ]r�B  (hh	e]r�B  (hj�)  e]r�B  (hh&e]r�B  (j�?  ]r�B  (hh	e]r�B  (hh	eeee]r�B  (hhee]r�B  (h]r�B  (hh e]r�B  (hh	e]r�B  (hhe]r�B  (h%h&eee]r�B  (j�=  ]r�B  (j�=  ]r�B  (j�=  ]r�B  (hj�)  e]r�B  (hj�)  e]r�B  (hjN  e]r�B  (j�=  ]r�B  (hh	e]r�B  (hj�)  e]r�B  (hh&e]r�B  (j�?  ]r�B  (hh	e]r�B  (hh	eeee]r�B  (hhee]r�B  (h]r�B  (hh e]r�B  (hh	e]r�B  (hhe]r�B  (h%h&eeej�B  j�B  j�B  j�B  ]r�B  (j�=  ]r�B  (j�=  ]r�B  (j�=  ]r�B  (hj�)  e]r�B  (hj�)  e]r�B  (hjN  e]r�B  (j�=  ]r�B  (hh	e]r�B  (hj�)  e]r�B  (hh&e]r�B  (j�?  ]r�B  (hh	e]r�B  (hh	eeee]r�B  (hhee]r�B  (h]r�B  (hh e]r�B  (hh	e]r�B  (hhe]r�B  (h%h&eeej�B  j�B  j�B  j�B  j�B  j�B  j�B  ]r�B  (j�=  ]r�B  (j�=  ]r C  (j�=  ]rC  (hj�)  e]rC  (hh	e]rC  (hjN  e]rC  (j�=  ]rC  (hh	e]rC  (hj�)  e]rC  (hh&e]rC  (j�?  ]r	C  (hh	e]r
C  (hh	eeee]rC  (hhee]rC  (h]rC  (hh e]rC  (hh	e]rC  (hhe]rC  (h%h&eeej�B  j�B  j�B  j�B  j�B  j�B  j�B  ]rC  (j�=  ]rC  (j�=  ]rC  (j�=  ]rC  (hj�)  e]rC  (hh	e]rC  (hjN  e]rC  (j�=  ]rC  (hj�)  e]rC  (hj�)  e]rC  (hh&e]rC  (j�?  ]rC  (hh	e]rC  (hh	eeee]rC  (hhee]rC  (h]r C  (hh e]r!C  (hh	e]r"C  (hhe]r#C  (h%h&eeejC  jC  jC  jC  jC  jC  jC  jC  jC  jC  ]r$C  (j�=  ]r%C  (j�=  ]r&C  (j�=  ]r'C  (hj�)  e]r(C  (hh	e]r)C  (hjN  e]r*C  (j�=  ]r+C  (hj�)  e]r,C  (hj�)  e]r-C  (hh&e]r.C  (j�?  ]r/C  (hh	e]r0C  (hh	eeee]r1C  (hhee]r2C  (h]r3C  (hh e]r4C  (hh	e]r5C  (hhe]r6C  (h%h&eee]r7C  (j�=  ]r8C  (j�=  ]r9C  (j�=  ]r:C  (hj�)  e]r;C  (hh	e]r<C  (hjN  e]r=C  (j�=  ]r>C  (hj�)  e]r?C  (hj�)  e]r@C  (hh&e]rAC  (j�?  ]rBC  (hh	e]rCC  (hh	eeee]rDC  (hhee]rEC  (h]rFC  (hh e]rGC  (hh	e]rHC  (hhe]rIC  (h%h&eee]rJC  (j�=  ]rKC  (j�=  ]rLC  (j�=  ]rMC  (hj�)  e]rNC  (hj�)  e]rOC  (hjN  e]rPC  (j�=  ]rQC  (hj�)  e]rRC  (hj�)  e]rSC  (hh&e]rTC  (j�?  ]rUC  (hh	e]rVC  (hh	eeee]rWC  (hhee]rXC  (h]rYC  (hh e]rZC  (hh	e]r[C  (hhe]r\C  (h%h&eeejJC  jJC  ]r]C  (j�=  ]r^C  (j�=  ]r_C  (j�=  ]r`C  (hj�)  e]raC  (hj�)  e]rbC  (hjN  e]rcC  (j�=  ]rdC  (hj�)  e]reC  (hj�)  e]rfC  (hh&e]rgC  (j�?  ]rhC  (hh	e]riC  (hh	eeee]rjC  (hhee]rkC  (h]rlC  (hh e]rmC  (hh	e]rnC  (hhe]roC  (h%h&eeej]C  j]C  j]C  j]C  j]C  j]C  j]C  j]C  ]rpC  (j�=  ]rqC  (j�=  ]rrC  (j�=  ]rsC  (hj�)  e]rtC  (hj�)  e]ruC  (hjN  e]rvC  (j�=  ]rwC  (hj�)  e]rxC  (hj�)  e]ryC  (hh&e]rzC  (j�?  ]r{C  (hh	e]r|C  (hh	eeee]r}C  (hhee]r~C  (h]rC  (hh e]r�C  (hh	e]r�C  (hhe]r�C  (h%h&eeejpC  ]r�C  (j�=  ]r�C  (j�=  ]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hj�)  e]r�C  (hjN  e]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hj�)  e]r�C  (hh&e]r�C  (j�?  ]r�C  (hh	e]r�C  (hh	eeee]r�C  (hhee]r�C  (h]r�C  (hh e]r�C  (hh	e]r�C  (hhe]r�C  (h%h&eeej�C  ]r�C  (j�=  ]r�C  (j�=  ]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hj�)  e]r�C  (hjN  e]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hh	e]r�C  (hh&e]r�C  (j�?  ]r�C  (hh	e]r�C  (hh	eeee]r�C  (hhee]r�C  (h]r�C  (hh e]r�C  (hh	e]r�C  (hhe]r�C  (h%h&eeej�C  j�C  j�C  ]r�C  (j�=  ]r�C  (j�=  ]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hj�)  e]r�C  (hjN  e]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hh	e]r�C  (hh&e]r�C  (j�?  ]r�C  (hh	e]r�C  (hh	eeee]r�C  (hhee]r�C  (h]r�C  (hh e]r�C  (hh	e]r�C  (hhe]r�C  (h%h&eee]r�C  (j�=  ]r�C  (j�=  ]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hj�)  e]r�C  (hjN  e]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hj�)  e]r�C  (hh&e]r�C  (j�?  ]r�C  (hh	e]r�C  (hh	eeee]r�C  (hhee]r�C  (h]r�C  (hh e]r�C  (hh	e]r�C  (hhe]r�C  (h%h&eee]r�C  (j�=  ]r�C  (j�=  ]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hh	e]r�C  (hjN  e]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hj�)  e]r�C  (hh&e]r�C  (j�?  ]r�C  (hh	e]r�C  (hh	eeee]r�C  (hhee]r�C  (h]r�C  (hh e]r�C  (hh	e]r�C  (hhe]r�C  (h%h&eee]r�C  (j�=  ]r�C  (j�=  ]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hh	e]r�C  (hjN  e]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hj�)  e]r�C  (hh&e]r�C  (j�?  ]r�C  (hh	e]r�C  (hh	eeee]r�C  (hhee]r�C  (h]r�C  (hh e]r�C  (hh	e]r�C  (hhe]r�C  (h%h&eeej�C  j�C  j�C  ]r�C  (j�=  ]r�C  (j�=  ]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hh	e]r�C  (hjN  e]r�C  (j�=  ]r�C  (hj�)  e]r�C  (hj�)  e]r�C  (hh&e]r�C  (j�?  ]r D  (hh	e]rD  (hh	eeee]rD  (hhee]rD  (h]rD  (hh e]rD  (hh	e]rD  (hhe]rD  (h%h&eee]rD  (j�=  ]r	D  (j�=  ]r
D  (j�=  ]rD  (hj�)  e]rD  (hh	e]rD  (hjN  e]rD  (j�=  ]rD  (hj�)  e]rD  (hj�)  e]rD  (hh&e]rD  (j�?  ]rD  (hh	e]rD  (hh	eeee]rD  (hhee]rD  (h]rD  (hh e]rD  (hh	e]rD  (hhe]rD  (h%h&eeejD  jD  ]rD  (j�=  ]rD  (j�=  ]rD  (j�=  ]rD  (hj�)  e]rD  (hh	e]r D  (hjN  e]r!D  (j�=  ]r"D  (hj�)  e]r#D  (hj�)  e]r$D  (hh&e]r%D  (j�?  ]r&D  (hh	e]r'D  (hh	eeee]r(D  (hhee]r)D  (h]r*D  (hh e]r+D  (hh	e]r,D  (hhe]r-D  (h%h&eee]r.D  (j�=  ]r/D  (j�=  ]r0D  (j�=  ]r1D  (hj�)  e]r2D  (hh	e]r3D  (hjN  e]r4D  (j�=  ]r5D  (hj�)  e]r6D  (hj�)  e]r7D  (hh&e]r8D  (j�?  ]r9D  (hh	e]r:D  (hh	eeee]r;D  (hhee]r<D  (h]r=D  (hh e]r>D  (hh	e]r?D  (hhe]r@D  (h%h&eeej.D  ]rAD  (j�=  ]rBD  (j�=  ]rCD  (j�=  ]rDD  (hj�)  e]rED  (hj�)  e]rFD  (hjN  e]rGD  (j�=  ]rHD  (hj�)  e]rID  (hj�)  e]rJD  (hh&e]rKD  (j�?  ]rLD  (hh	e]rMD  (hh	eeee]rND  (hhee]rOD  (h]rPD  (hh e]rQD  (hh	e]rRD  (hhe]rSD  (h%h&eeejAD  jAD  jAD  ]rTD  (j�=  ]rUD  (j�=  ]rVD  (j�=  ]rWD  (hj�)  e]rXD  (hj�)  e]rYD  (hjN  e]rZD  (j�=  ]r[D  (hj�)  e]r\D  (hj�)  e]r]D  (hh&e]r^D  (j�?  ]r_D  (hh	e]r`D  (hh	eeee]raD  (hhee]rbD  (h]rcD  (hh e]rdD  (hh	e]reD  (hhe]rfD  (h%h&eeejTD  jTD  jTD  ]rgD  (j�=  ]rhD  (j�=  ]riD  (j�=  ]rjD  (hj�)  e]rkD  (hj�)  e]rlD  (hjN  e]rmD  (j�=  ]rnD  (hj�)  e]roD  (hj�)  e]rpD  (hh&e]rqD  (j�?  ]rrD  (hh	e]rsD  (hh	eeee]rtD  (hhee]ruD  (h]rvD  (hh e]rwD  (hh	e]rxD  (hhe]ryD  (h%h&eeejgD  ]rzD  (j�=  ]r{D  (j�=  ]r|D  (j�=  ]r}D  (hj�)  e]r~D  (hj�)  e]rD  (hjN  e]r�D  (j�=  ]r�D  (hj�)  e]r�D  (hj�)  e]r�D  (hh&e]r�D  (j�?  ]r�D  (hh	e]r�D  (hh	eeee]r�D  (hhee]r�D  (h]r�D  (hh e]r�D  (hh	e]r�D  (hhe]r�D  (h%h&eee]r�D  (j�=  ]r�D  (j�=  ]r�D  (j�=  ]r�D  (hj�)  e]r�D  (hj�)  e]r�D  (hjN  e]r�D  (j�=  ]r�D  (hj�)  e]r�D  (hj�)  e]r�D  (hh&e]r�D  (j�?  ]r�D  (hh	e]r�D  (hh	eeee]r�D  (hhee]r�D  (h]r�D  (hh e]r�D  (hh	e]r�D  (hhe]r�D  (h%h&eeej�D  j�D  j�D  j�D  j�D  ]r�D  (j�=  ]r�D  (j�=  ]r�D  (j�=  ]r�D  (hj�)  e]r�D  (hj�)  e]r�D  (hjN  e]r�D  (j�=  ]r�D  (hh	e]r�D  (hj�)  e]r�D  (hh&e]r�D  (j�?  ]r�D  (hh	e]r�D  (hh	eeee]r�D  (hhee]r�D  (h]r�D  (hh e]r�D  (hh	e]r�D  (hhe]r�D  (h%h&eeej�D  j�D  j�D  ]r�D  (j�=  ]r�D  (j�=  ]r�D  (j�=  ]r�D  (hj�)  e]r�D  (hj�)  e]r�D  (hjN  e]r�D  (j�=  ]r�D  (hh	e]r�D  (hj�)  e]r�D  (hh&e]r�D  (j�?  ]r�D  (hh	e]r�D  (hh	eeee]r�D  (hhee]r�D  (h]r�D  (hh e]r�D  (hh	e]r�D  (hhe]r�D  (h%h&eeej�D  ]r�D  (j�=  ]r�D  (j�=  ]r�D  (j�=  ]r�D  (hj�)  e]r�D  (hj�)  e]r�D  (hjN  e]r�D  (j�=  ]r�D  (hh	e]r�D  (hj�)  e]r�D  (hh&e]r�D  (j�?  ]r�D  (hh	e]r�D  (hh	eeee]r�D  (hhee]r�D  (h]r�D  (hh e]r�D  (hh	e]r�D  (hhe]r�D  (h%h&eee]r�D  (j�=  ]r�D  (j�=  ]r�D  (j�=  ]r�D  (hj�)  e]r�D  (hj�)  e]r�D  (hjN  e]r�D  (j�=  ]r�D  (hh	e]r�D  (hj�)  e]r�D  (hh&e]r�D  (j�?  ]r�D  (hh	e]r�D  (hh	eeee]r�D  (hhee]r�D  (h]r�D  (hh e]r�D  (hh	e]r�D  (hhe]r�D  (h%h&eeej�D  j�D  j�D  ]r�D  (j�=  ]r�D  (j�=  ]r�D  (j�=  ]r�D  (hj�)  e]r�D  (hj�)  e]r�D  (hjN  e]r�D  (j�=  ]r�D  (hh	e]r�D  (hj�)  e]r�D  (hh&e]r�D  (j�?  ]r�D  (hh	e]r�D  (hh	eeee]r�D  (hhee]r�D  (h]r�D  (hh e]r�D  (hh	e]r�D  (hhe]r�D  (h%h&eeej�D  j�D  j�D  j�D  j�D  j�D  j�D  ]r�D  (j�=  ]r E  (j�=  ]rE  (j�=  ]rE  (hj�)  e]rE  (hj�)  e]rE  (hjN  e]rE  (j�=  ]rE  (hh	e]rE  (hj�)  e]rE  (hh&e]r	E  (j�?  ]r
E  (hh	e]rE  (hh	eeee]rE  (hhee]rE  (h]rE  (hh e]rE  (hh	e]rE  (hhe]rE  (h%h&eeej�D  ]rE  (j�=  ]rE  (j�=  ]rE  (j�=  ]rE  (hj�)  e]rE  (hj�)  e]rE  (hjN  e]rE  (j�=  ]rE  (hh	e]rE  (hj�)  e]rE  (hh&e]rE  (j�?  ]rE  (hh	e]rE  (hh	eeee]rE  (hhee]r E  (h]r!E  (hh e]r"E  (hh	e]r#E  (hhe]r$E  (h%h&eee]r%E  (j�=  ]r&E  (j�=  ]r'E  (j�=  ]r(E  (hj�)  e]r)E  (hj�)  e]r*E  (hjN  e]r+E  (j�=  ]r,E  (hh	e]r-E  (hj�)  e]r.E  (hh&e]r/E  (j�?  ]r0E  (hh	e]r1E  (hh	eeee]r2E  (hhee]r3E  (h]r4E  (hh e]r5E  (hh	e]r6E  (hhe]r7E  (h%h&eeej%E  j%E  j%E  ]r8E  (j�=  ]r9E  (j�=  ]r:E  (j�=  ]r;E  (hj�)  e]r<E  (hj�)  e]r=E  (hjN  e]r>E  (j�=  ]r?E  (hh	e]r@E  (hj�)  e]rAE  (hh&e]rBE  (j�?  ]rCE  (hh	e]rDE  (hh	eeee]rEE  (hhee]rFE  (h]rGE  (hh e]rHE  (hh	e]rIE  (hhe]rJE  (h%h&eeej8E  ]rKE  (j�=  ]rLE  (j�=  ]rME  (j�=  ]rNE  (hj�)  e]rOE  (hj�)  e]rPE  (hjN  e]rQE  (j�=  ]rRE  (hh	e]rSE  (hj�)  e]rTE  (hh&e]rUE  (j�?  ]rVE  (hh	e]rWE  (hh	eeee]rXE  (hhee]rYE  (h]rZE  (hh e]r[E  (hh	e]r\E  (hhe]r]E  (h%h&eee]r^E  (j�=  ]r_E  (j�=  ]r`E  (j�=  ]raE  (hh	e]rbE  (hj�)  e]rcE  (hjN  e]rdE  (j�=  ]reE  (hh	e]rfE  (hj�)  e]rgE  (hh&e]rhE  (j�?  ]riE  (hh	e]rjE  (hh	eeee]rkE  (hhee]rlE  (h]rmE  (hh e]rnE  (hh	e]roE  (hhe]rpE  (h%h&eee]rqE  (j�=  ]rrE  (j�=  ]rsE  (j�=  ]rtE  (hh	e]ruE  (hj�)  e]rvE  (hjN  e]rwE  (j�=  ]rxE  (hj�)  e]ryE  (hj�)  e]rzE  (hh&e]r{E  (j�?  ]r|E  (hh	e]r}E  (hh	eeee]r~E  (hhee]rE  (h]r�E  (hh e]r�E  (hh	e]r�E  (hhe]r�E  (h%h&eeejqE  jqE  jqE  jqE  ]r�E  (j�=  ]r�E  (j�=  ]r�E  (j�=  ]r�E  (hh	e]r�E  (hj�)  e]r�E  (hjN  e]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hh&e]r�E  (j�?  ]r�E  (hh	e]r�E  (hh	eeee]r�E  (hhee]r�E  (h]r�E  (hh e]r�E  (hh	e]r�E  (hhe]r�E  (h%h&eee]r�E  (j�=  ]r�E  (j�=  ]r�E  (j�=  ]r�E  (hh	e]r�E  (hj�)  e]r�E  (hjN  e]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hh&e]r�E  (j�?  ]r�E  (hh	e]r�E  (hh	eeee]r�E  (hhee]r�E  (h]r�E  (hh e]r�E  (hh	e]r�E  (hhe]r�E  (h%h&eeej�E  ]r�E  (j�=  ]r�E  (j�=  ]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hjN  e]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hh&e]r�E  (j�?  ]r�E  (hh	e]r�E  (hh	eeee]r�E  (hhee]r�E  (h]r�E  (hh e]r�E  (hh	e]r�E  (hhe]r�E  (h%h&eee]r�E  (j�=  ]r�E  (j�=  ]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hjN  e]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hh&e]r�E  (j�?  ]r�E  (hh	e]r�E  (hh	eeee]r�E  (hhee]r�E  (h]r�E  (hh e]r�E  (hh	e]r�E  (hhe]r�E  (h%h&eeej�E  j�E  j�E  j�E  j�E  j�E  j�E  j�E  j�E  ]r�E  (j�=  ]r�E  (j�=  ]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hjN  e]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hh&e]r�E  (j�?  ]r�E  (hh	e]r�E  (hh	eeee]r�E  (hhee]r�E  (h]r�E  (hh e]r�E  (hh	e]r�E  (hhe]r�E  (h%h&eeej�E  ]r�E  (j�=  ]r�E  (j�=  ]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hjN  e]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hh&e]r�E  (j�?  ]r�E  (hh	e]r�E  (hh	eeee]r�E  (hhee]r�E  (h]r�E  (hh e]r�E  (hh	e]r�E  (hhe]r�E  (h%h&eee]r�E  (j�=  ]r�E  (j�=  ]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hjN  e]r�E  (j�=  ]r�E  (hj�)  e]r�E  (hj�)  e]r�E  (hh&e]r F  (j�?  ]rF  (hh	e]rF  (hh	eeee]rF  (hhee]rF  (h]rF  (hh e]rF  (hh	e]rF  (hhe]rF  (h%h&eeej�E  j�E  ]r	F  (j�=  ]r
F  (j�=  ]rF  (j�=  ]rF  (hj�)  e]rF  (hj�)  e]rF  (hjN  e]rF  (j�=  ]rF  (hj�)  e]rF  (hj�)  e]rF  (hh&e]rF  (j�?  ]rF  (hh	e]rF  (hh	eeee]rF  (hhee]rF  (h]rF  (hh e]rF  (hh	e]rF  (hhe]rF  (h%h&eeej	F  j	F  j	F  ]rF  (j�=  ]rF  (j�=  ]rF  (j�=  ]rF  (hj�)  e]r F  (hj�)  e]r!F  (hjN  e]r"F  (j�=  ]r#F  (hj�)  e]r$F  (hj�)  e]r%F  (hh&e]r&F  (j�?  ]r'F  (hh	e]r(F  (hh	eeee]r)F  (hhee]r*F  (h]r+F  (hh e]r,F  (hh	e]r-F  (hhe]r.F  (h%h&eee]r/F  (j�=  ]r0F  (j�=  ]r1F  (j�=  ]r2F  (hj�)  e]r3F  (hj�)  e]r4F  (hjN  e]r5F  (j�=  ]r6F  (hj�)  e]r7F  (hj�)  e]r8F  (hh&e]r9F  (j�?  ]r:F  (hh	e]r;F  (hh	eeee]r<F  (hhee]r=F  (h]r>F  (hh e]r?F  (hh	e]r@F  (hhe]rAF  (h%h&eeej/F  j/F  j/F  j/F  j/F  j/F  j/F  j/F  j/F  ]rBF  (j�=  ]rCF  (j�=  ]rDF  (j�=  ]rEF  (hj�)  e]rFF  (hj�)  e]rGF  (hjN  e]rHF  (j�=  ]rIF  (hj�)  e]rJF  (hj�)  e]rKF  (hh&e]rLF  (j�?  ]rMF  (hh	e]rNF  (hh	eeee]rOF  (hhee]rPF  (h]rQF  (hh e]rRF  (hh	e]rSF  (hhe]rTF  (h%h&eee]rUF  (j�=  ]rVF  (j�=  ]rWF  (j�=  ]rXF  (hj�)  e]rYF  (hj�)  e]rZF  (hjN  e]r[F  (j�=  ]r\F  (hj�)  e]r]F  (hj�)  e]r^F  (hh&e]r_F  (j�?  ]r`F  (hh	e]raF  (hh	eeee]rbF  (hhee]rcF  (h]rdF  (hh e]reF  (hh	e]rfF  (hhe]rgF  (h%h&eee]rhF  (j�=  ]riF  (j�=  ]rjF  (j�=  ]rkF  (hj�)  e]rlF  (hj�)  e]rmF  (hjN  e]rnF  (j�=  ]roF  (hj�)  e]rpF  (hj�)  e]rqF  (hh&e]rrF  (X	   Next-MoversF  ]rtF  (hh	e]ruF  (hh	eeee]rvF  (hhee]rwF  (h]rxF  (hh e]ryF  (hh	e]rzF  (hhe]r{F  (h%h&eee]r|F  (j�=  ]r}F  (j�=  ]r~F  (j�=  ]rF  (hj�)  e]r�F  (hj�)  e]r�F  (hjN  e]r�F  (j�=  ]r�F  (hj�)  e]r�F  (hj�)  e]r�F  (hh&e]r�F  (jsF  ]r�F  (hh	e]r�F  (hh	eeee]r�F  (hhee]r�F  (h]r�F  (hh e]r�F  (hh	e]r�F  (hhe]r�F  (h%h&eeej|F  j|F  j|F  j|F  j|F  j|F  ]r�F  (j�=  ]r�F  (j�=  ]r�F  (j�=  ]r�F  (hj�)  e]r�F  (hj�)  e]r�F  (hjN  e]r�F  (j�=  ]r�F  (hh	e]r�F  (hj�)  e]r�F  (hh&e]r�F  (jsF  ]r�F  (hh	e]r�F  (hh	eeee]r�F  (hhee]r�F  (h]r�F  (hh e]r�F  (hh	e]r�F  (hhe]r�F  (h%h&eee]r�F  (j�=  ]r�F  (j�=  ]r�F  (j�=  ]r�F  (hj�)  e]r�F  (hj�)  e]r�F  (hjN  e]r�F  (j�=  ]r�F  (hh	e]r�F  (hj�)  e]r�F  (hh&e]r�F  (jsF  ]r�F  (hh	e]r�F  (hh	eeee]r�F  (hhee]r�F  (h]r�F  (hh e]r�F  (hh	e]r�F  (hhe]r�F  (h%h&eeej�F  j�F  j�F  j�F  j�F  ]r�F  (j�=  ]r�F  (j�=  ]r�F  (j�=  ]r�F  (hj�)  e]r�F  (hj�)  e]r�F  (hjN  e]r�F  (j�=  ]r�F  (hh	e]r�F  (hj�)  e]r�F  (hh&e]r�F  (jsF  ]r�F  (hh	e]r�F  (hh	eeee]r�F  (hhee]r�F  (h]r�F  (hh e]r�F  (hh	e]r�F  (hhe]r�F  (h%h&eeej�F  ]r�F  (j�=  ]r�F  (j�=  ]r�F  (j�=  ]r�F  (hj�)  e]r�F  (hj�)  e]r�F  (hjN  e]r�F  (j�=  ]r�F  (hh	e]r�F  (hj�)  e]r�F  (hh&e]r�F  (X	   Next-Mover�F  ]r�F  (hh	e]r�F  (hh	eeee]r�F  (hhee]r�F  (h]r�F  (hh e]r�F  (hh	e]r�F  (hhe]r�F  (h%h&eee]r�F  (j�=  ]r�F  (j�=  ]r�F  (j�=  ]r�F  (hj�)  e]r�F  (hj�)  e]r�F  (hjN  e]r�F  (j�=  ]r�F  (hh	e]r�F  (hj�)  e]r�F  (hh&e]r�F  (j�F  ]r�F  (hh	e]r�F  (hh	eeee]r�F  (hhee]r�F  (h]r�F  (hh e]r�F  (hh	e]r�F  (hhe]r�F  (h%h&eeej�F  ]r�F  (j�=  ]r�F  (j�=  ]r�F  (j�=  ]r�F  (hj�)  e]r�F  (hj�)  e]r�F  (hjN  e]r�F  (j�=  ]r�F  (hj�)  e]r�F  (hj�)  e]r�F  (hh&e]r�F  (j�F  ]r�F  (hh	e]r�F  (hh	eeee]r�F  (hhee]r�F  (h]r�F  (hh e]r�F  (hh	e]r G  (hhe]rG  (h%h&eee]rG  (j�=  ]rG  (j�=  ]rG  (j�=  ]rG  (hj�)  e]rG  (hj�)  e]rG  (hjN  e]rG  (j�=  ]r	G  (hh	e]r
G  (hj�)  e]rG  (hh&e]rG  (j�F  ]rG  (hh	e]rG  (hh	eeee]rG  (hhee]rG  (h]rG  (hh e]rG  (hh	e]rG  (hhe]rG  (h%h&eeejG  ]rG  (j�=  ]rG  (j�=  ]rG  (j�=  ]rG  (hj�)  e]rG  (hj�)  e]rG  (hjN  e]rG  (j�=  ]rG  (hh	e]rG  (hj�)  e]rG  (hh&e]rG  (j�F  ]r G  (hh	e]r!G  (hh	eeee]r"G  (hhee]r#G  (h]r$G  (hh e]r%G  (hh	e]r&G  (hhe]r'G  (h%h&eee]r(G  (j�=  ]r)G  (j�=  ]r*G  (j�=  ]r+G  (hj�)  e]r,G  (hj�)  e]r-G  (hjN  e]r.G  (j�=  ]r/G  (hh	e]r0G  (hj�)  e]r1G  (hh&e]r2G  (j�F  ]r3G  (hh	e]r4G  (hh	eeee]r5G  (hhee]r6G  (h]r7G  (hh e]r8G  (hh	e]r9G  (hhe]r:G  (h%h&eee]r;G  (j�=  ]r<G  (j�=  ]r=G  (j�=  ]r>G  (hj�)  e]r?G  (hj�)  e]r@G  (hjN  e]rAG  (j�=  ]rBG  (hh	e]rCG  (hj�)  e]rDG  (hh&e]rEG  (j�F  ]rFG  (hh	e]rGG  (hh	eeee]rHG  (hhee]rIG  (h]rJG  (hh e]rKG  (hh	e]rLG  (hhe]rMG  (h%h&eeej;G  j;G  ]rNG  (j�=  ]rOG  (j�=  ]rPG  (j�=  ]rQG  (hj�)  e]rRG  (hj�)  e]rSG  (hjN  e]rTG  (j�=  ]rUG  (hh	e]rVG  (hj�)  e]rWG  (hh&e]rXG  (j�F  ]rYG  (hh	e]rZG  (hh	eeee]r[G  (hhee]r\G  (h]r]G  (hh e]r^G  (hh	e]r_G  (hhe]r`G  (h%h&eee]raG  (j�=  ]rbG  (j�=  ]rcG  (j�=  ]rdG  (hj�)  e]reG  (hj�)  e]rfG  (hjN  e]rgG  (j�=  ]rhG  (hh	e]riG  (hj�)  e]rjG  (hh&e]rkG  (j�F  ]rlG  (hh	e]rmG  (hh	eeee]rnG  (hhee]roG  (h]rpG  (hh e]rqG  (hh	e]rrG  (hhe]rsG  (h%h&eeejaG  jaG  jaG  ]rtG  (j�=  ]ruG  (j�=  ]rvG  (j�=  ]rwG  (hh	e]rxG  (hj�)  e]ryG  (hjN  e]rzG  (j�=  ]r{G  (hh	e]r|G  (hj�)  e]r}G  (hh&e]r~G  (j�F  ]rG  (hh	e]r�G  (hh	eeee]r�G  (hhee]r�G  (h]r�G  (hh e]r�G  (hh	e]r�G  (hhe]r�G  (h%h&eeejtG  jtG  jtG  jtG  jtG  jtG  jtG  jtG  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hjN  e]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hh&e]r�G  (j�F  ]r�G  (hh	e]r�G  (hh	eeee]r�G  (hhee]r�G  (h]r�G  (hh e]r�G  (hh	e]r�G  (hhe]r�G  (h%h&eeej�G  j�G  j�G  j�G  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hjN  e]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hh&e]r�G  (j�F  ]r�G  (hh	e]r�G  (hh	eeee]r�G  (hhee]r�G  (h]r�G  (hh e]r�G  (hh	e]r�G  (hhe]r�G  (h%h&eeej�G  j�G  j�G  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hjN  e]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hh&e]r�G  (j�F  ]r�G  (hh	e]r�G  (hh	eeee]r�G  (hhee]r�G  (h]r�G  (hh e]r�G  (hh	e]r�G  (hhe]r�G  (h%h&eeej�G  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hjN  e]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hh&e]r�G  (j�F  ]r�G  (hh	e]r�G  (hh	eeee]r�G  (hhee]r�G  (h]r�G  (hh e]r�G  (hh	e]r�G  (hhe]r�G  (h%h&eeej�G  j�G  j�G  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hjN  e]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hh&e]r�G  (j�F  ]r�G  (hh	e]r�G  (hh	eeee]r�G  (hhee]r�G  (h]r�G  (hh e]r�G  (hh	e]r�G  (hhe]r�G  (h%h&eee]r�G  (j�=  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hjN  e]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hh&e]r�G  (j�F  ]r�G  (hh	e]r�G  (hh	eeee]r�G  (hhee]r�G  (h]r�G  (hh e]r�G  (hh	e]r�G  (hhe]r�G  (h%h&eeej�G  j�G  j�G  j�G  j�G  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (j�=  ]r�G  (hh	e]r�G  (hj�)  e]r�G  (hjN  e]r�G  (j�=  ]r H  (hh	e]rH  (hj�)  e]rH  (hh&e]rH  (j�F  ]rH  (hh	e]rH  (hh	eeee]rH  (hhee]rH  (h]rH  (hh e]r	H  (hh	e]r
H  (hhe]rH  (h%h&eeej�G  ]rH  (j�=  ]rH  (j�=  ]rH  (j�=  ]rH  (hh	e]rH  (hj�)  e]rH  (hjN  e]rH  (j�=  ]rH  (hh	e]rH  (hj�)  e]rH  (hh&e]rH  (j�F  ]rH  (hh	e]rH  (hh	eeee]rH  (hhee]rH  (h]rH  (hh e]rH  (hh	e]rH  (hhe]rH  (h%h&eeejH  jH  jH  jH  jH  jH  ]rH  (j�=  ]r H  (j�=  ]r!H  (j�=  ]r"H  (hh	e]r#H  (hj�)  e]r$H  (hjN  e]r%H  (j�=  ]r&H  (hh	e]r'H  (hj�)  e]r(H  (hh&e]r)H  (j�F  ]r*H  (hh	e]r+H  (hh	eeee]r,H  (hhee]r-H  (h]r.H  (hh e]r/H  (hh	e]r0H  (hhe]r1H  (h%h&eeejH  jH  jH  jH  jH  jH  jH  jH  jH  ]r2H  (j�=  ]r3H  (j�=  ]r4H  (j�=  ]r5H  (hh	e]r6H  (hj�)  e]r7H  (hjN  e]r8H  (j�=  ]r9H  (hh	e]r:H  (hj�)  e]r;H  (hh&e]r<H  (j�F  ]r=H  (hh	e]r>H  (hh	eeee]r?H  (hhee]r@H  (h]rAH  (hh e]rBH  (hh	e]rCH  (hhe]rDH  (h%h&eeej2H  j2H  j2H  j2H  j2H  j2H  j2H  j2H  j2H  ]rEH  (j�=  ]rFH  (j�=  ]rGH  (j�=  ]rHH  (hh	e]rIH  (hj�)  e]rJH  (hjN  e]rKH  (j�=  ]rLH  (hh	e]rMH  (hj�)  e]rNH  (hh&e]rOH  (j�F  ]rPH  (hh	e]rQH  (hh	eeee]rRH  (hhee]rSH  (h]rTH  (hh e]rUH  (hh	e]rVH  (hhe]rWH  (h%h&eeejEH  jEH  ]rXH  (j�=  ]rYH  (j�=  ]rZH  (j�=  ]r[H  (hh	e]r\H  (hj�)  e]r]H  (hjN  e]r^H  (j�=  ]r_H  (hh	e]r`H  (hj�)  e]raH  (hh&e]rbH  (j�F  ]rcH  (hh	e]rdH  (hh	eeee]reH  (hhee]rfH  (h]rgH  (hh e]rhH  (hh	e]riH  (hhe]rjH  (h%h&eeejXH  ]rkH  (j�=  ]rlH  (j�=  ]rmH  (j�=  ]rnH  (hh	e]roH  (hj�)  e]rpH  (hjN  e]rqH  (j�=  ]rrH  (hh	e]rsH  (hj�)  e]rtH  (hh&e]ruH  (j�F  ]rvH  (hh	e]rwH  (hh	eeee]rxH  (hhee]ryH  (h]rzH  (hh e]r{H  (hh	e]r|H  (hhe]r}H  (h%h&eeejkH  jkH  jkH  jkH  jkH  jkH  jkH  jkH  ]r~H  (j�=  ]rH  (j�=  ]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hjN  e]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hh&e]r�H  (j�F  ]r�H  (hh	e]r�H  (hh	eeee]r�H  (hhee]r�H  (h]r�H  (hh e]r�H  (hh	e]r�H  (hhe]r�H  (h%h&eeej~H  j~H  j~H  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hjN  e]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hh&e]r�H  (j�F  ]r�H  (hh	e]r�H  (hh	eeee]r�H  (hhee]r�H  (h]r�H  (hh e]r�H  (hh	e]r�H  (hhe]r�H  (h%h&eeej�H  j�H  j�H  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hjN  e]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hh&e]r�H  (j�F  ]r�H  (hh	e]r�H  (hh	eeee]r�H  (hhee]r�H  (h]r�H  (hh e]r�H  (hh	e]r�H  (hhe]r�H  (h%h&eeej�H  j�H  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hjN  e]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hh&e]r�H  (j�F  ]r�H  (hh	e]r�H  (hh	eeee]r�H  (hhee]r�H  (h]r�H  (hh e]r�H  (hh	e]r�H  (hhe]r�H  (h%h&eeej�H  j�H  j�H  j�H  j�H  j�H  j�H  j�H  j�H  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hjN  e]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hh&e]r�H  (j�F  ]r�H  (hh	e]r�H  (hh	eeee]r�H  (hhee]r�H  (h]r�H  (hh e]r�H  (hh	e]r�H  (hhe]r�H  (h%h&eeej�H  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hjN  e]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hh&e]r�H  (j�F  ]r�H  (hh	e]r�H  (hh	eeee]r�H  (hhee]r�H  (h]r�H  (hh e]r�H  (hh	e]r�H  (hhe]r�H  (h%h&eeej�H  j�H  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (j�=  ]r�H  (hh	e]r�H  (hj�)  e]r�H  (hjN  e]r�H  (j�=  ]r�H  (hj�)  e]r�H  (hj�)  e]r�H  (hh&e]r�H  (j�F  ]r�H  (hh	e]r�H  (hh	eeee]r�H  (hhee]r�H  (h]r�H  (hh e]r I  (hh	e]rI  (hhe]rI  (h%h&eeej�H  j�H  j�H  ]rI  (j�=  ]rI  (j�=  ]rI  (j�=  ]rI  (hh	e]rI  (hj�)  e]rI  (hjN  e]r	I  (j�=  ]r
I  (hj�)  e]rI  (hj�)  e]rI  (hh&e]rI  (j�F  ]rI  (hh	e]rI  (hh	eeee]rI  (hhee]rI  (h]rI  (hh e]rI  (hh	e]rI  (hhe]rI  (h%h&eeejI  ]rI  (j�=  ]rI  (j�=  ]rI  (j�=  ]rI  (hh	e]rI  (hj�)  e]rI  (hjN  e]rI  (j�=  ]rI  (hj�)  e]rI  (hj�)  e]rI  (hh&e]r I  (j�F  ]r!I  (hh	e]r"I  (hh	eeee]r#I  (hhee]r$I  (h]r%I  (hh e]r&I  (hh	e]r'I  (hhe]r(I  (h%h&eeejI  jI  jI  jI  jI  jI  jI  jI  ]r)I  (j�=  ]r*I  (j�=  ]r+I  (j�=  ]r,I  (hh	e]r-I  (hj�)  e]r.I  (hjN  e]r/I  (j�=  ]r0I  (hj�)  e]r1I  (hh	e]r2I  (hh&e]r3I  (j�F  ]r4I  (hh	e]r5I  (hh	eeee]r6I  (hhee]r7I  (h]r8I  (hh e]r9I  (hh	e]r:I  (hhe]r;I  (h%h&eeej)I  j)I  j)I  j)I  j)I  ]r<I  (j�=  ]r=I  (j�=  ]r>I  (j�=  ]r?I  (hh	e]r@I  (hj�)  e]rAI  (hjN  e]rBI  (j�=  ]rCI  (hj�)  e]rDI  (hh	e]rEI  (hh&e]rFI  (j�F  ]rGI  (hh	e]rHI  (hh	eeee]rII  (hhee]rJI  (h]rKI  (hh e]rLI  (hh	e]rMI  (hhe]rNI  (h%h&eeej<I  j<I  j<I  j<I  j<I  j<I  j<I  j<I  ]rOI  (j�=  ]rPI  (j�=  ]rQI  (j�=  ]rRI  (hh	e]rSI  (hj�)  e]rTI  (hjN  e]rUI  (j�=  ]rVI  (hj�)  e]rWI  (hh	e]rXI  (hh&e]rYI  (j�F  ]rZI  (hh	e]r[I  (hh	eeee]r\I  (hhee]r]I  (h]r^I  (hh e]r_I  (hh	e]r`I  (hhe]raI  (h%h&eeejOI  jOI  jOI  jOI  ]rbI  (j�=  ]rcI  (j�=  ]rdI  (j�=  ]reI  (hh	e]rfI  (hj�)  e]rgI  (hjN  e]rhI  (j�=  ]riI  (hj�)  e]rjI  (hj�)  e]rkI  (hh&e]rlI  (j�F  ]rmI  (hh	e]rnI  (hh	eeee]roI  (hhee]rpI  (h]rqI  (hh e]rrI  (hh	e]rsI  (hhe]rtI  (h%h&eee]ruI  (j�=  ]rvI  (j�=  ]rwI  (j�=  ]rxI  (hh	e]ryI  (hj�)  e]rzI  (hjN  e]r{I  (j�=  ]r|I  (hj�)  e]r}I  (hj�)  e]r~I  (hh&e]rI  (j�F  ]r�I  (hh	e]r�I  (hh	eeee]r�I  (hhee]r�I  (h]r�I  (hh e]r�I  (hh	e]r�I  (hhe]r�I  (h%h&eee]r�I  (j�=  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (hh	e]r�I  (hj�)  e]r�I  (hjN  e]r�I  (j�=  ]r�I  (hj�)  e]r�I  (hj�)  e]r�I  (hh&e]r�I  (j�F  ]r�I  (hh	e]r�I  (hh	eeee]r�I  (hhee]r�I  (h]r�I  (hh e]r�I  (hh	e]r�I  (hhe]r�I  (h%h&eeej�I  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (hh	e]r�I  (hj�)  e]r�I  (hjN  e]r�I  (j�=  ]r�I  (hj�)  e]r�I  (hj�)  e]r�I  (hh&e]r�I  (j�F  ]r�I  (hh	e]r�I  (hh	eeee]r�I  (hhee]r�I  (h]r�I  (hh e]r�I  (hh	e]r�I  (hhe]r�I  (h%h&eeej�I  j�I  j�I  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (hh	e]r�I  (hj�)  e]r�I  (hjN  e]r�I  (j�=  ]r�I  (hj�)  e]r�I  (hj�)  e]r�I  (hh&e]r�I  (j�F  ]r�I  (hh	e]r�I  (hh	eeee]r�I  (hhee]r�I  (h]r�I  (hh e]r�I  (hh	e]r�I  (hhe]r�I  (h%h&eeej�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (hh	e]r�I  (hj�)  e]r�I  (hjN  e]r�I  (j�=  ]r�I  (hj�)  e]r�I  (hj�)  e]r�I  (hh&e]r�I  (j�F  ]r�I  (hh	e]r�I  (hh	eeee]r�I  (hhee]r�I  (h]r�I  (hh e]r�I  (hh	e]r�I  (hhe]r�I  (h%h&eeej�I  j�I  j�I  j�I  j�I  j�I  j�I  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (hh	e]r�I  (hj�)  e]r�I  (hjN  e]r�I  (j�=  ]r�I  (hj�)  e]r�I  (hj�)  e]r�I  (hh&e]r�I  (j�F  ]r�I  (hh	e]r�I  (hh	eeee]r�I  (hhee]r�I  (h]r�I  (hh e]r�I  (hh	e]r�I  (hhe]r�I  (h%h&eeej�I  j�I  j�I  j�I  j�I  j�I  j�I  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (hh	e]r�I  (hj�)  e]r�I  (hjN  e]r�I  (j�=  ]r�I  (hj�)  e]r�I  (hj�)  e]r�I  (hh&e]r�I  (j�F  ]r�I  (hh	e]r�I  (hh	eeee]r�I  (hhee]r�I  (h]r�I  (hh e]r�I  (hh	e]r�I  (hhe]r�I  (h%h&eeej�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (j�=  ]r�I  (hh	e]r�I  (hj�)  e]r�I  (hjN  e]r J  (j�=  ]rJ  (hj�)  e]rJ  (hj�)  e]rJ  (hh&e]rJ  (j�F  ]rJ  (hh	e]rJ  (hh	eeee]rJ  (hhee]rJ  (h]r	J  (hh e]r
J  (hh	e]rJ  (hhe]rJ  (h%h&eeej�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  j�I  ]rJ  (j�=  ]rJ  (j�=  ]rJ  (j�=  ]rJ  (hh	e]rJ  (hj�)  e]rJ  (hjN  e]rJ  (j�=  ]rJ  (hj�)  e]rJ  (hh	e]rJ  (hh&e]rJ  (j�F  ]rJ  (hh	e]rJ  (hh	eeee]rJ  (hhee]rJ  (h]rJ  (hh e]rJ  (hh	e]rJ  (hhe]rJ  (h%h&eeejJ  jJ  jJ  jJ  jJ  jJ  jJ  jJ  ]r J  (j�=  ]r!J  (j�=  ]r"J  (j�=  ]r#J  (hh	e]r$J  (hj�)  e]r%J  (hjN  e]r&J  (j�=  ]r'J  (hj�)  e]r(J  (hh	e]r)J  (hh&e]r*J  (j�F  ]r+J  (hh	e]r,J  (hh	eeee]r-J  (hhee]r.J  (h]r/J  (hh e]r0J  (hh	e]r1J  (hhe]r2J  (h%h&eeej J  j J  j J  j J  ]r3J  (j�=  ]r4J  (j�=  ]r5J  (j�=  ]r6J  (hh	e]r7J  (hj�)  e]r8J  (hjN  e]r9J  (j�=  ]r:J  (hj�)  e]r;J  (hh	e]r<J  (hh&e]r=J  (j�F  ]r>J  (hh	e]r?J  (hh	eeee]r@J  (hhee]rAJ  (h]rBJ  (hh e]rCJ  (hh	e]rDJ  (hhe]rEJ  (h%h&eee]rFJ  (j�=  ]rGJ  (j�=  ]rHJ  (j�=  ]rIJ  (hh	e]rJJ  (hj�)  e]rKJ  (hjN  e]rLJ  (j�=  ]rMJ  (hj�)  e]rNJ  (hh	e]rOJ  (hh&e]rPJ  (j�F  ]rQJ  (hh	e]rRJ  (hh	eeee]rSJ  (hhee]rTJ  (h]rUJ  (hh e]rVJ  (hh	e]rWJ  (hhe]rXJ  (h%h&eee]rYJ  (j�=  ]rZJ  (j�=  ]r[J  (j�=  ]r\J  (hh	e]r]J  (hj�)  e]r^J  (hjN  e]r_J  (j�=  ]r`J  (hj�)  e]raJ  (hh	e]rbJ  (hh&e]rcJ  (j�F  ]rdJ  (hh	e]reJ  (hh	eeee]rfJ  (hhee]rgJ  (h]rhJ  (hh e]riJ  (hh	e]rjJ  (hhe]rkJ  (h%h&eeejYJ  jYJ  jYJ  jYJ  jYJ  ]rlJ  (j�=  ]rmJ  (j�=  ]rnJ  (j�=  ]roJ  (hh	e]rpJ  (hj�)  e]rqJ  (hjN  e]rrJ  (j�=  ]rsJ  (hj�)  e]rtJ  (hh	e]ruJ  (hh&e]rvJ  (j�F  ]rwJ  (hh	e]rxJ  (hh	eeee]ryJ  (hhee]rzJ  (h]r{J  (hh e]r|J  (hh	e]r}J  (hhe]r~J  (h%h&eeejlJ  jlJ  jlJ  ]rJ  (j�=  ]r�J  (j�=  ]r�J  (j�=  ]r�J  (hh	e]r�J  (hj�)  e]r�J  (hjN  e]r�J  (j�=  ]r�J  (hj�)  e]r�J  (hh	e]r�J  (hh&e]r�J  (X	   Next-Mover�J  ]r�J  (hh	e]r�J  (hh	eeee]r�J  (hhee]r�J  (h]r�J  (hh e]r�J  (hh	e]r�J  (hhe]r�J  (h%h&eee]r�J  (j�=  ]r�J  (j�=  ]r�J  (j�=  ]r�J  (hh	e]r�J  (hj�)  e]r�J  (hjN  e]r�J  (j�=  ]r�J  (hj�)  e]r�J  (hh	e]r�J  (hh&e]r�J  (j�J  ]r�J  (hh	e]r�J  (hh	eeee]r�J  (hhee]r�J  (h]r�J  (hh e]r�J  (hh	e]r�J  (hhe]r�J  (h%h&eeej�J  ]r�J  (j�=  ]r�J  (j�=  ]r�J  (j�=  ]r�J  (hh	e]r�J  (hj�)  e]r�J  (hjN  e]r�J  (j�=  ]r�J  (hj�)  e]r�J  (hh	e]r�J  (hh&e]r�J  (j�J  ]r�J  (hh	e]r�J  (hh	eeee]r�J  (hhee]r�J  (h]r�J  (hh e]r�J  (hh	e]r�J  (hhe]r�J  (h%h&eeej�J  j�J  j�J  j�J  j�J  j�J  j�J  ]r�J  (j�=  ]r�J  (j�=  ]r�J  (j�=  ]r�J  (hh	e]r�J  (hj�)  e]r�J  (hjN  e]r�J  (j�=  ]r�J  (hj�)  e]r�J  (hh	e]r�J  (hh&e]r�J  (j�J  ]r�J  (hh	e]r�J  (hh	eeee]r�J  (hhee]r�J  (h]r�J  (hh e]r�J  (hh	e]r�J  (hhe]r�J  (h%h&eeej�J  ]r�J  (j�=  ]r�J  (j�=  ]r�J  (j�=  ]r�J  (hh	e]r�J  (hj�)  e]r�J  (hjN  e]r�J  (j�=  ]r�J  (hj�)  e]r�J  (hh	e]r�J  (hh&e]r�J  (j�J  ]r�J  (hh	e]r�J  (hh	eeee]r�J  (hhee]r�J  (h]r�J  (hh e]r�J  (hh	e]r�J  (hhe]r�J  (h%h&eee]r�J  (j�=  ]r�J  (j�=  ]r�J  (j�=  ]r�J  (hh	e]r�J  (hj�)  e]r�J  (hjN  e]r�J  (j�=  ]r�J  (hj�)  e]r�J  (hh	e]r�J  (hh&e]r�J  (j�J  ]r�J  (hh	e]r�J  (hh	eeee]r�J  (hhee]r�J  (h]r�J  (hh e]r�J  (hh	e]r�J  (hhe]r�J  (h%h&eee]r�J  (j�=  ]r�J  (j�=  ]r�J  (j�=  ]r�J  (hh	e]r�J  (hj�)  e]r�J  (hjN  e]r�J  (j�=  ]r�J  (hj�)  e]r�J  (hh	e]r�J  (hh&e]r�J  (j�J  ]r�J  (hh	e]r�J  (hh	eeee]r�J  (hhee]r K  (h]rK  (hh e]rK  (hh	e]rK  (hhe]rK  (h%h&eeej�J  ]rK  (j�=  ]rK  (j�=  ]rK  (j�=  ]rK  (hh	e]r	K  (hj�)  e]r
K  (hjN  e]rK  (j�=  ]rK  (hj�)  e]rK  (hh	e]rK  (hh&e]rK  (j�J  ]rK  (hh	e]rK  (hh	eeee]rK  (hhee]rK  (h]rK  (hh e]rK  (hh	e]rK  (hhe]rK  (h%h&eeejK  jK  ]rK  (j�=  ]rK  (j�=  ]rK  (j�=  ]rK  (hh	e]rK  (hj�)  e]rK  (hjN  e]rK  (j�=  ]rK  (hj�)  e]r K  (hh	e]r!K  (hh&e]r"K  (j�J  ]r#K  (hh	e]r$K  (hh	eeee]r%K  (hhee]r&K  (h]r'K  (hh e]r(K  (hh	e]r)K  (hhe]r*K  (h%h&eeejK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  jK  ]r+K  (j�=  ]r,K  (j�=  ]r-K  (j�=  ]r.K  (hh	e]r/K  (hj�)  e]r0K  (hjN  e]r1K  (j�=  ]r2K  (hj�)  e]r3K  (hh	e]r4K  (hh&e]r5K  (j�J  ]r6K  (hh	e]r7K  (hh	eeee]r8K  (hhee]r9K  (h]r:K  (hh e]r;K  (hh	e]r<K  (hhe]r=K  (h%h&eeej+K  j+K  j+K  ]r>K  (j�=  ]r?K  (j�=  ]r@K  (j�=  ]rAK  (hh	e]rBK  (hj�)  e]rCK  (hjN  e]rDK  (j�=  ]rEK  (hj�)  e]rFK  (hh	e]rGK  (hh&e]rHK  (j�J  ]rIK  (hh	e]rJK  (hh	eeee]rKK  (hhee]rLK  (h]rMK  (hh e]rNK  (hh	e]rOK  (hhe]rPK  (h%h&eeej>K  ]rQK  (j�=  ]rRK  (j�=  ]rSK  (j�=  ]rTK  (hh	e]rUK  (hj�)  e]rVK  (hjN  e]rWK  (j�=  ]rXK  (hj�)  e]rYK  (hh	e]rZK  (hh&e]r[K  (j�J  ]r\K  (hh	e]r]K  (hh	eeee]r^K  (hhee]r_K  (h]r`K  (hh e]raK  (hh	e]rbK  (hhe]rcK  (h%h&eeejQK  ]rdK  (j�=  ]reK  (j�=  ]rfK  (j�=  ]rgK  (hh	e]rhK  (hj�)  e]riK  (hjN  e]rjK  (j�=  ]rkK  (hj�)  e]rlK  (hh	e]rmK  (hh&e]rnK  (j�J  ]roK  (hh	e]rpK  (hh	eeee]rqK  (hhee]rrK  (h]rsK  (hh e]rtK  (hh	e]ruK  (hhe]rvK  (h%h&eee]rwK  (j�=  ]rxK  (j�=  ]ryK  (j�=  ]rzK  (hh	e]r{K  (hj�)  e]r|K  (hjN  e]r}K  (j�=  ]r~K  (hj�)  e]rK  (hh	e]r�K  (hh&e]r�K  (j�J  ]r�K  (hh	e]r�K  (hh	eeee]r�K  (hhee]r�K  (h]r�K  (hh e]r�K  (hh	e]r�K  (hhe]r�K  (h%h&eeejwK  ]r�K  (j�=  ]r�K  (j�=  ]r�K  (j�=  ]r�K  (hh	e]r�K  (hj�)  e]r�K  (hjN  e]r�K  (j�=  ]r�K  (hj�)  e]r�K  (hh	e]r�K  (hh&e]r�K  (j�J  ]r�K  (hh	e]r�K  (hh	eeee]r�K  (hhee]r�K  (h]r�K  (hh e]r�K  (hh	e]r�K  (hhe]r�K  (h%h&eeej�K  j�K  j�K  j�K  j�K  j�K  ]r�K  (j�=  ]r�K  (j�=  ]r�K  (j�=  ]r�K  (hh	e]r�K  (hj�)  e]r�K  (hjN  e]r�K  (j�=  ]r�K  (hj�)  e]r�K  (hh	e]r�K  (hh&e]r�K  (j�J  ]r�K  (hh	e]r�K  (hh	eeee]r�K  (hhee]r�K  (h]r�K  (hh e]r�K  (hh	e]r�K  (hhe]r�K  (h%h&eee]r�K  (j�=  ]r�K  (j�=  ]r�K  (j�=  ]r�K  (hh	e]r�K  (hj�)  e]r�K  (hjN  e]r�K  (j�=  ]r�K  (hj�)  e]r�K  (hh	e]r�K  (hh&e]r�K  (j�J  ]r�K  (hh	e]r�K  (hh	eeee]r�K  (hhee]r�K  (h]r�K  (hh e]r�K  (hh	e]r�K  (hhe]r�K  (h%h&eeej�K  j�K  j�K  j�K  j�K  j�K  ]r�K  (j�=  ]r�K  (j�=  ]r�K  (j�=  ]r�K  (hh	e]r�K  (hj�)  e]r�K  (hjN  e]r�K  (j�=  ]r�K  (hj�)  e]r�K  (hh	e]r�K  (hh&e]r�K  (j�J  ]r�K  (hh	e]r�K  (hh	eeee]r�K  (hhee]r�K  (h]r�K  (hh e]r�K  (hh	e]r�K  (hhe]r�K  (h%h&eee]r�K  (j�=  ]r�K  (j�=  ]r�K  (j�=  ]r�K  (hh	e]r�K  (hj�)  e]r�K  (hjN  e]r�K  (j�=  ]r�K  (hj�)  e]r�K  (hh	e]r�K  (hh&e]r�K  (j�J  ]r�K  (hh	e]r�K  (hh	eeee]r�K  (hhee]r�K  (h]r�K  (hh e]r�K  (hh	e]r�K  (hhe]r�K  (h%h&eeej�K  j�K  j�K  j�K  j�K  j�K  j�K  ]r�K  (j�=  ]r�K  (j�=  ]r�K  (j�=  ]r�K  (hh	e]r�K  (hj�)  e]r�K  (hjN  e]r�K  (j�=  ]r�K  (hj�)  e]r�K  (hh	e]r�K  (hh&e]r�K  (j�J  ]r�K  (hh	e]r�K  (hh	eeee]r�K  (hhee]r�K  (h]r�K  (hh e]r�K  (hh	e]r�K  (hhe]r�K  (h%h&eee]r�K  (j�=  ]r�K  (j�=  ]r�K  (j�=  ]r�K  (hh	e]r L  (hj�)  e]rL  (hjN  e]rL  (j�=  ]rL  (hj�)  e]rL  (hj�)  e]rL  (hh&e]rL  (j�J  ]rL  (hh	e]rL  (hh	eeee]r	L  (hhee]r
L  (h]rL  (hh e]rL  (hh	e]rL  (hhe]rL  (h%h&eeej�K  j�K  j�K  j�K  j�K  j�K  j�K  ]rL  (j�=  ]rL  (j�=  ]rL  (j�=  ]rL  (hh	e]rL  (hj�)  e]rL  (hjN  e]rL  (j�=  ]rL  (hh	e]rL  (hj�)  e]rL  (hh&e]rL  (j�J  ]rL  (hh	e]rL  (hh	eeee]rL  (hhee]rL  (h]rL  (hh e]rL  (hh	e]r L  (hhe]r!L  (h%h&eeejL  ]r"L  (j�=  ]r#L  (j�=  ]r$L  (j�=  ]r%L  (hh	e]r&L  (hj�)  e]r'L  (hjN  e]r(L  (j�=  ]r)L  (hh	e]r*L  (hj�)  e]r+L  (hh&e]r,L  (j�J  ]r-L  (hh	e]r.L  (hh	eeee]r/L  (hhee]r0L  (h]r1L  (hh e]r2L  (hh	e]r3L  (hhe]r4L  (h%h&eeej"L  j"L  j"L  j"L  j"L  j"L  ]r5L  (j�=  ]r6L  (j�=  ]r7L  (j�=  ]r8L  (hh	e]r9L  (hj�)  e]r:L  (hjN  e]r;L  (j�=  ]r<L  (hh	e]r=L  (hj�)  e]r>L  (hh&e]r?L  (j�J  ]r@L  (hh	e]rAL  (hh	eeee]rBL  (hhee]rCL  (h]rDL  (hh e]rEL  (hh	e]rFL  (hhe]rGL  (h%h&eee]rHL  (j�=  ]rIL  (j�=  ]rJL  (j�=  ]rKL  (hh	e]rLL  (hj�)  e]rML  (hjN  e]rNL  (j�=  ]rOL  (hh	e]rPL  (hj�)  e]rQL  (hh&e]rRL  (j�J  ]rSL  (hh	e]rTL  (hh	eeee]rUL  (hhee]rVL  (h]rWL  (hh e]rXL  (hh	e]rYL  (hhe]rZL  (h%h&eeejHL  jHL  jHL  ]r[L  (j�=  ]r\L  (j�=  ]r]L  (j�=  ]r^L  (hh	e]r_L  (hj�)  e]r`L  (hjN  e]raL  (j�=  ]rbL  (hh	e]rcL  (hj�)  e]rdL  (hh&e]reL  (j�J  ]rfL  (hh	e]rgL  (hh	eeee]rhL  (hhee]riL  (h]rjL  (hh e]rkL  (hh	e]rlL  (hhe]rmL  (h%h&eeej[L  j[L  j[L  ]rnL  (j�=  ]roL  (j�=  ]rpL  (j�=  ]rqL  (hh	e]rrL  (hj�)  e]rsL  (hjN  e]rtL  (j�=  ]ruL  (hh	e]rvL  (hj�)  e]rwL  (hh&e]rxL  (j�J  ]ryL  (hh	e]rzL  (hh	eeee]r{L  (hhee]r|L  (h]r}L  (hh e]r~L  (hh	e]rL  (hhe]r�L  (h%h&eeejnL  jnL  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hjN  e]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hh&e]r�L  (j�J  ]r�L  (hh	e]r�L  (hh	eeee]r�L  (hhee]r�L  (h]r�L  (hh e]r�L  (hh	e]r�L  (hhe]r�L  (h%h&eeej�L  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hjN  e]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hh&e]r�L  (j�J  ]r�L  (hh	e]r�L  (hh	eeee]r�L  (hhee]r�L  (h]r�L  (hh e]r�L  (hh	e]r�L  (hhe]r�L  (h%h&eeej�L  j�L  j�L  j�L  j�L  j�L  j�L  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hjN  e]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hh&e]r�L  (j�J  ]r�L  (hh	e]r�L  (hh	eeee]r�L  (hhee]r�L  (h]r�L  (hh e]r�L  (hh	e]r�L  (hhe]r�L  (h%h&eeej�L  j�L  j�L  j�L  j�L  j�L  j�L  j�L  j�L  j�L  j�L  j�L  j�L  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hjN  e]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hh&e]r�L  (j�J  ]r�L  (hh	e]r�L  (hh	eeee]r�L  (hhee]r�L  (h]r�L  (hh e]r�L  (hh	e]r�L  (hhe]r�L  (h%h&eeej�L  j�L  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hjN  e]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hh&e]r�L  (j�J  ]r�L  (hh	e]r�L  (hh	eeee]r�L  (hhee]r�L  (h]r�L  (hh e]r�L  (hh	e]r�L  (hhe]r�L  (h%h&eeej�L  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hjN  e]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hh&e]r�L  (j�J  ]r�L  (hh	e]r�L  (hh	eeee]r�L  (hhee]r�L  (h]r�L  (hh e]r�L  (hh	e]r�L  (hhe]r�L  (h%h&eee]r�L  (j�=  ]r�L  (j�=  ]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hjN  e]r�L  (j�=  ]r�L  (hh	e]r�L  (hj�)  e]r�L  (hh&e]r�L  (j�J  ]r�L  (hh	e]r�L  (hh	eeee]r M  (hhee]rM  (h]rM  (hh e]rM  (hh	e]rM  (hhe]rM  (h%h&eee]rM  (j�=  ]rM  (j�=  ]rM  (j�=  ]r	M  (hh	e]r
M  (hj�)  e]rM  (hjN  e]rM  (j�=  ]rM  (hh	e]rM  (hj�)  e]rM  (hh&e]rM  (j�J  ]rM  (hh	e]rM  (hh	eeee]rM  (hhee]rM  (h]rM  (hh e]rM  (hh	e]rM  (hhe]rM  (h%h&eeejM  jM  ]rM  (j�=  ]rM  (j�=  ]rM  (j�=  ]rM  (hh	e]rM  (hj�)  e]rM  (hjN  e]rM  (j�=  ]r M  (hj�)  e]r!M  (hj�)  e]r"M  (hh&e]r#M  (j�J  ]r$M  (hh	e]r%M  (hh	eeee]r&M  (hhee]r'M  (h]r(M  (hh e]r)M  (hh	e]r*M  (hhe]r+M  (h%h&eeejM  jM  jM  jM  jM  jM  ]r,M  (j�=  ]r-M  (j�=  ]r.M  (j�=  ]r/M  (hh	e]r0M  (hj�)  e]r1M  (hjN  e]r2M  (j�=  ]r3M  (hj�)  e]r4M  (hj�)  e]r5M  (hh&e]r6M  (j�J  ]r7M  (hh	e]r8M  (hh	eeee]r9M  (hhee]r:M  (h]r;M  (hh e]r<M  (hh	e]r=M  (hhe]r>M  (h%h&eee]r?M  (j�=  ]r@M  (j�=  ]rAM  (j�=  ]rBM  (hh	e]rCM  (hj�)  e]rDM  (hjN  e]rEM  (j�=  ]rFM  (hj�)  e]rGM  (hj�)  e]rHM  (hh&e]rIM  (j�J  ]rJM  (hh	e]rKM  (hh	eeee]rLM  (hhee]rMM  (h]rNM  (hh e]rOM  (hh	e]rPM  (hhe]rQM  (h%h&eeej?M  j?M  j?M  j?M  j?M  j?M  j?M  ]rRM  (j�=  ]rSM  (j�=  ]rTM  (j�=  ]rUM  (hh	e]rVM  (hj�)  e]rWM  (hjN  e]rXM  (j�=  ]rYM  (hj�)  e]rZM  (hj�)  e]r[M  (hh&e]r\M  (X	   Next-Mover]M  ]r^M  (hh	e]r_M  (hh	eeee]r`M  (hhee]raM  (h]rbM  (hh e]rcM  (hh	e]rdM  (hhe]reM  (h%h&eeejRM  jRM  jRM  jRM  jRM  ]rfM  (j�=  ]rgM  (j�=  ]rhM  (j�=  ]riM  (hh	e]rjM  (hj�)  e]rkM  (hjN  e]rlM  (j�=  ]rmM  (hj�)  e]rnM  (hj�)  e]roM  (hh&e]rpM  (j]M  ]rqM  (hh	e]rrM  (hh	eeee]rsM  (hhee]rtM  (h]ruM  (hh e]rvM  (hh	e]rwM  (hhe]rxM  (h%h&eeejfM  jfM  jfM  jfM  jfM  jfM  jfM  jfM  jfM  jfM  jfM  ]ryM  (j�=  ]rzM  (j�=  ]r{M  (j�=  ]r|M  (hh	e]r}M  (hj�)  e]r~M  (hjN  e]rM  (j�=  ]r�M  (hj�)  e]r�M  (hj�)  e]r�M  (hh&e]r�M  (j]M  ]r�M  (hh	e]r�M  (hh	eeee]r�M  (hhee]r�M  (h]r�M  (hh e]r�M  (hh	e]r�M  (hhe]r�M  (h%h&eeejyM  ]r�M  (j�=  ]r�M  (j�=  ]r�M  (j�=  ]r�M  (hh	e]r�M  (hj�)  e]r�M  (hjN  e]r�M  (j�=  ]r�M  (hj�)  e]r�M  (hj�)  e]r�M  (hh&e]r�M  (j]M  ]r�M  (hh	e]r�M  (hh	eeee]r�M  (hhee]r�M  (h]r�M  (hh e]r�M  (hh	e]r�M  (hhe]r�M  (h%h&eeej�M  ]r�M  (j�=  ]r�M  (j�=  ]r�M  (j�=  ]r�M  (hh	e]r�M  (hj�)  e]r�M  (hjN  e]r�M  (j�=  ]r�M  (hj�)  e]r�M  (hj�)  e]r�M  (hh&e]r�M  (j]M  ]r�M  (hh	e]r�M  (hh	eeee]r�M  (hhee]r�M  (h]r�M  (hh e]r�M  (hh	e]r�M  (hhe]r�M  (h%h&eeej�M  j�M  ]r�M  (j�=  ]r�M  (j�=  ]r�M  (j�=  ]r�M  (hj�)  e]r�M  (hj�)  e]r�M  (hjN  e]r�M  (j�=  ]r�M  (hj�)  e]r�M  (hj�)  e]r�M  (hh&e]r�M  (j]M  ]r�M  (hh	e]r�M  (hh	eeee]r�M  (hhee]r�M  (h]r�M  (hh e]r�M  (hh	e]r�M  (hhe]r�M  (h%h&eee]r�M  (j�=  ]r�M  (j�=  ]r�M  (j�=  ]r�M  (hj�)  e]r�M  (hj�)  e]r�M  (hjN  e]r�M  (j�=  ]r�M  (hj�)  e]r�M  (hj�)  e]r�M  (hh&e]r�M  (j]M  ]r�M  (hh	e]r�M  (hh	eeee]r�M  (hhee]r�M  (h]r�M  (hh e]r�M  (hh	e]r�M  (hhe]r�M  (h%h&eeej�M  ]r�M  (j�=  ]r�M  (j�=  ]r�M  (j�=  ]r�M  (hj�)  e]r�M  (hj�)  e]r�M  (hjN  e]r�M  (j�=  ]r�M  (hj�)  e]r�M  (hj�)  e]r�M  (hh&e]r�M  (j]M  ]r�M  (hh	e]r�M  (hh	eeee]r�M  (hhee]r�M  (h]r�M  (hh e]r�M  (hh	e]r�M  (hhe]r�M  (h%h&eee]r�M  (j�=  ]r�M  (j�=  ]r�M  (j�=  ]r�M  (hj�)  e]r�M  (hj�)  e]r�M  (hjN  e]r�M  (j�=  ]r�M  (hj�)  e]r�M  (hj�)  e]r�M  (hh&e]r�M  (j]M  ]r�M  (hh	e]r�M  (hh	eeee]r�M  (hhee]r�M  (h]r�M  (hh e]r�M  (hh	e]r�M  (hhe]r�M  (h%h&eeej�M  j�M  ]r�M  (j�=  ]r�M  (j�=  ]r N  (j�=  ]rN  (hj�)  e]rN  (hj�)  e]rN  (hjN  e]rN  (j�=  ]rN  (hj�)  e]rN  (hj�)  e]rN  (hh&e]rN  (j]M  ]r	N  (hh	e]r
N  (hh	eeee]rN  (hhee]rN  (h]rN  (hh e]rN  (hh	e]rN  (hhe]rN  (h%h&eeej�M  j�M  ]rN  (j�=  ]rN  (j�=  ]rN  (j�=  ]rN  (hj�)  e]rN  (hj�)  e]rN  (hjN  e]rN  (j�=  ]rN  (hj�)  e]rN  (hj�)  e]rN  (hh&e]rN  (j]M  ]rN  (hh	e]rN  (hh	eeee]rN  (hhee]rN  (h]r N  (hh e]r!N  (hh	e]r"N  (hhe]r#N  (h%h&eeejN  jN  ]r$N  (j�=  ]r%N  (j�=  ]r&N  (j�=  ]r'N  (hj�)  e]r(N  (hj�)  e]r)N  (hjN  e]r*N  (j�=  ]r+N  (hj�)  e]r,N  (hj�)  e]r-N  (hh&e]r.N  (j]M  ]r/N  (hh	e]r0N  (hh	eeee]r1N  (hhee]r2N  (h]r3N  (hh e]r4N  (hh	e]r5N  (hhe]r6N  (h%h&eeej$N  j$N  j$N  j$N  ]r7N  (j�=  ]r8N  (j�=  ]r9N  (j�=  ]r:N  (hj�)  e]r;N  (hj�)  e]r<N  (hjN  e]r=N  (j�=  ]r>N  (hj�)  e]r?N  (hj�)  e]r@N  (hh&e]rAN  (j]M  ]rBN  (hh	e]rCN  (hh	eeee]rDN  (hhee]rEN  (h]rFN  (hh e]rGN  (hh	e]rHN  (hhe]rIN  (h%h&eeej7N  j7N  ]rJN  (j�=  ]rKN  (j�=  ]rLN  (j�=  ]rMN  (hj�)  e]rNN  (hj�)  e]rON  (hjN  e]rPN  (j�=  ]rQN  (hj�)  e]rRN  (hj�)  e]rSN  (hh&e]rTN  (j]M  ]rUN  (hh	e]rVN  (hh	eeee]rWN  (hhee]rXN  (h]rYN  (hh e]rZN  (hh	e]r[N  (hhe]r\N  (h%h&eeejJN  jJN  ]r]N  (j�=  ]r^N  (j�=  ]r_N  (j�=  ]r`N  (hj�)  e]raN  (hj�)  e]rbN  (hjN  e]rcN  (j�=  ]rdN  (hj�)  e]reN  (hj�)  e]rfN  (hh&e]rgN  (j]M  ]rhN  (hh	e]riN  (hh	eeee]rjN  (hhee]rkN  (h]rlN  (hh e]rmN  (hh	e]rnN  (hhe]roN  (h%h&eeej]N  j]N  j]N  j]N  ]rpN  (j�=  ]rqN  (j�=  ]rrN  (j�=  ]rsN  (hj�)  e]rtN  (hj�)  e]ruN  (hjN  e]rvN  (j�=  ]rwN  (hj�)  e]rxN  (hj�)  e]ryN  (hh&e]rzN  (j]M  ]r{N  (hh	e]r|N  (hh	eeee]r}N  (hhee]r~N  (h]rN  (hh e]r�N  (hh	e]r�N  (hhe]r�N  (h%h&eeejpN  jpN  jpN  jpN  jpN  jpN  jpN  jpN  jpN  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hj�)  e]r�N  (hjN  e]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hj�)  e]r�N  (hh&e]r�N  (j]M  ]r�N  (hh	e]r�N  (hh	eeee]r�N  (hhee]r�N  (h]r�N  (hh e]r�N  (hh	e]r�N  (hhe]r�N  (h%h&eeej�N  j�N  j�N  j�N  j�N  j�N  j�N  j�N  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hj�)  e]r�N  (hjN  e]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hj�)  e]r�N  (hh&e]r�N  (j]M  ]r�N  (hh	e]r�N  (hh	eeee]r�N  (hhee]r�N  (h]r�N  (hh e]r�N  (hh	e]r�N  (hhe]r�N  (h%h&eee]r�N  (j�=  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hh	e]r�N  (hjN  e]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hj�)  e]r�N  (hh&e]r�N  (j]M  ]r�N  (hh	e]r�N  (hh	eeee]r�N  (hhee]r�N  (h]r�N  (hh e]r�N  (hh	e]r�N  (hhe]r�N  (h%h&eeej�N  j�N  j�N  j�N  j�N  j�N  j�N  j�N  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hh	e]r�N  (hjN  e]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hj�)  e]r�N  (hh&e]r�N  (j]M  ]r�N  (hh	e]r�N  (hh	eeee]r�N  (hhee]r�N  (h]r�N  (hh e]r�N  (hh	e]r�N  (hhe]r�N  (h%h&eeej�N  j�N  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hh	e]r�N  (hjN  e]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hj�)  e]r�N  (hh&e]r�N  (j]M  ]r�N  (hh	e]r�N  (hh	eeee]r�N  (hhee]r�N  (h]r�N  (hh e]r�N  (hh	e]r�N  (hhe]r�N  (h%h&eeej�N  j�N  j�N  j�N  j�N  j�N  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hh	e]r�N  (hjN  e]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hj�)  e]r�N  (hh&e]r�N  (j]M  ]r�N  (hh	e]r�N  (hh	eeee]r�N  (hhee]r�N  (h]r�N  (hh e]r�N  (hh	e]r�N  (hhe]r�N  (h%h&eeej�N  j�N  j�N  j�N  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hh	e]r�N  (hjN  e]r�N  (j�=  ]r�N  (hj�)  e]r�N  (hj�)  e]r�N  (hh&e]r�N  (j]M  ]r O  (hh	e]rO  (hh	eeee]rO  (hhee]rO  (h]rO  (hh e]rO  (hh	e]rO  (hhe]rO  (h%h&eeej�N  j�N  j�N  j�N  j�N  j�N  j�N  j�N  j�N  ]rO  (j�=  ]r	O  (j�=  ]r
O  (j�=  ]rO  (hj�)  e]rO  (hh	e]rO  (hjN  e]rO  (j�=  ]rO  (hj�)  e]rO  (hj�)  e]rO  (hh&e]rO  (j]M  ]rO  (hh	e]rO  (hh	eeee]rO  (hhee]rO  (h]rO  (hh e]rO  (hh	e]rO  (hhe]rO  (h%h&eeejO  jO  jO  jO  jO  jO  jO  jO  jO  jO  jO  jO  jO  jO  jO  ]rO  (j�=  ]rO  (j�=  ]rO  (j�=  ]rO  (hj�)  e]rO  (hh	e]r O  (hjN  e]r!O  (j�=  ]r"O  (hj�)  e]r#O  (hj�)  e]r$O  (hh&e]r%O  (j]M  ]r&O  (hh	e]r'O  (hh	eeee]r(O  (hhee]r)O  (h]r*O  (hh e]r+O  (hh	e]r,O  (hhe]r-O  (h%h&eeejO  jO  jO  jO  ]r.O  (j�=  ]r/O  (j�=  ]r0O  (j�=  ]r1O  (hj�)  e]r2O  (hh	e]r3O  (hjN  e]r4O  (j�=  ]r5O  (hj�)  e]r6O  (hj�)  e]r7O  (hh&e]r8O  (j]M  ]r9O  (hh	e]r:O  (hh	eeee]r;O  (hhee]r<O  (h]r=O  (hh e]r>O  (hh	e]r?O  (hhe]r@O  (h%h&eeej.O  j.O  ]rAO  (j�=  ]rBO  (j�=  ]rCO  (j�=  ]rDO  (hj�)  e]rEO  (hh	e]rFO  (hjN  e]rGO  (j�=  ]rHO  (hj�)  e]rIO  (hj�)  e]rJO  (hh&e]rKO  (j]M  ]rLO  (hh	e]rMO  (hh	eeee]rNO  (hhee]rOO  (h]rPO  (hh e]rQO  (hh	e]rRO  (hhe]rSO  (h%h&eee]rTO  (j�=  ]rUO  (j�=  ]rVO  (j�=  ]rWO  (hj�)  e]rXO  (hh	e]rYO  (hjN  e]rZO  (j�=  ]r[O  (hj�)  e]r\O  (hj�)  e]r]O  (hh&e]r^O  (j]M  ]r_O  (hh	e]r`O  (hh	eeee]raO  (hhee]rbO  (h]rcO  (hh e]rdO  (hh	e]reO  (hhe]rfO  (h%h&eee]rgO  (j�=  ]rhO  (j�=  ]riO  (j�=  ]rjO  (hj�)  e]rkO  (hh	e]rlO  (hjN  e]rmO  (j�=  ]rnO  (hj�)  e]roO  (hj�)  e]rpO  (hh&e]rqO  (j]M  ]rrO  (hh	e]rsO  (hh	eeee]rtO  (hhee]ruO  (h]rvO  (hh e]rwO  (hh	e]rxO  (hhe]ryO  (h%h&eee]rzO  (j�=  ]r{O  (j�=  ]r|O  (j�=  ]r}O  (hj�)  e]r~O  (hh	e]rO  (hjN  e]r�O  (j�=  ]r�O  (hj�)  e]r�O  (hj�)  e]r�O  (hh&e]r�O  (j]M  ]r�O  (hh	e]r�O  (hh	eeee]r�O  (hhee]r�O  (h]r�O  (hh e]r�O  (hh	e]r�O  (hhe]r�O  (h%h&eee]r�O  (j�=  ]r�O  (j�=  ]r�O  (j�=  ]r�O  (hj�)  e]r�O  (hh	e]r�O  (hjN  e]r�O  (j�=  ]r�O  (hh	e]r�O  (hj�)  e]r�O  (hh&e]r�O  (j]M  ]r�O  (hh	e]r�O  (hh	eeee]r�O  (hhee]r�O  (h]r�O  (hh e]r�O  (hh	e]r�O  (hhe]r�O  (h%h&eeej�O  j�O  j�O  j�O  ]r�O  (j�=  ]r�O  (j�=  ]r�O  (j�=  ]r�O  (hj�)  e]r�O  (hh	e]r�O  (hjN  e]r�O  (j�=  ]r�O  (hh	e]r�O  (hj�)  e]r�O  (hh&e]r�O  (j]M  ]r�O  (hh	e]r�O  (hh	eeee]r�O  (hhee]r�O  (h]r�O  (hh e]r�O  (hh	e]r�O  (hhe]r�O  (h%h&eeej�O  ]r�O  (j�=  ]r�O  (j�=  ]r�O  (j�=  ]r�O  (hj�)  e]r�O  (hh	e]r�O  (hjN  e]r�O  (j�=  ]r�O  (hh	e]r�O  (hj�)  e]r�O  (hh&e]r�O  (X	   Next-Mover�O  ]r�O  (hh	e]r�O  (hh	eeee]r�O  (hhee]r�O  (h]r�O  (hh e]r�O  (hh	e]r�O  (hhe]r�O  (h%h&eeej�O  ]r�O  (j�=  ]r�O  (j�=  ]r�O  (j�=  ]r�O  (hj�)  e]r�O  (hh	e]r�O  (hjN  e]r�O  (j�=  ]r�O  (hh	e]r�O  (hj�)  e]r�O  (hh&e]r�O  (j�O  ]r�O  (hh	e]r�O  (hh	eeee]r�O  (hhee]r�O  (h]r�O  (hh e]r�O  (hh	e]r�O  (hhe]r�O  (h%h&eeee.