�]q (X   pickupqK�qX   putdownqKK�q�qhK�qhKK�q�qhK%�q	hK%K�q
�qhK�qhKcnumpy.core.multiarray
scalar
qcnumpy
dtype
qX   i4qK K�qRq(KX   <qNNNJ����J����K tqbC   q�qRq�q�qhK�qhKhhC   q�qRq�q�qhK�qhKK�q �q!hK�q"hKK�q#�q$hK%�q%hK%K�q&�q'hK�q(hKhhC   q)�q*Rq+�q,�q-hK�q.hKhhC   q/�q0Rq1�q2�q3hK�q4hKhhC   q5�q6Rq7�q8�q9hK%�q:hK%K�q;�q<hK�q=hKhhC   q>�q?Rq@�qA�qBhK�qChKK�qD�qEhK�qFhKK�qG�qHhK%�qIhK%K�qJ�qKhK�qLhKhhC   qM�qNRqO�qP�qQhK�qRhKhhC   qS�qTRqU�qV�qWhK�qXhKK�qY�qZhK�q[hKK�q\�q]hK�q^hKK�q_�q`hK�qahKhhC   qb�qcRqd�qe�qfhK�qghKhhC   qh�qiRqj�qk�qlhK�qmhKK�qn�qohK%�qphK%K�qq�qrhK�qshKK�qt�quhK�qvhKhhC   qw�qxRqy�qz�q{hK�q|hKK�q}�q~hK%�qhK%K�q��q�hK�q�hKhhC   q��q�Rq��q��q�hK�q�hKhhC   q��q�Rq��q��q�hK�q�hKhhC   q��q�Rq��q��q�hK%�q�hK%K�q��q�hK�q�hKK�q��q�hK�q�hKK�q��q�hK�q�hKhhC   q��q�Rq��q��q�hK%�q�hK%K�q��q�hK�q�hKK�q��q�hK�q�hKhhC   q��q�Rq��q��q�hK�q�hKK�q��q�hK%�q�hK%K�q��q�hK�q�hKhhC   q��q�Rq��q��q�hK�q�hKhhC   q��q�Rq��q��q�hK�q�hKK�qq�hK�q�hKK�qņq�hK�q�hKK�qȆq�hK%�q�hK%K�qˆq�hK�q�hKhhC   qΆq�RqЇqцq�hK�q�hKK�qԆq�hK�q�hKhhC   q׆q�Rqهqچq�hK�q�hKhhC   q݆q�Rq߇q��q�hK%�q�hK%K�q�q�hK�q�hKK�q�q�hK�q�hKhhC   q�q�Rq�q�q�hK�q�hKK�q�q�hK�q�hKhhC   q�q�Rq�q��q�hK�q�hKhhC   q��q�Rq��q��q�hK�q�hKK�q��q�hK%�r   hK%K�r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr	  �r
  �r  hK�r  hKK�r  �r  hK�r  hKK�r  �r  hK%�r  hK%K�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK%�r  hK%K�r  �r  hK�r  hKhhC   r  �r   Rr!  �r"  �r#  hK�r$  hKK�r%  �r&  hK�r'  hKhhC   r(  �r)  Rr*  �r+  �r,  hK�r-  hKK�r.  �r/  hK�r0  hKK�r1  �r2  hK�r3  hKhhC   r4  �r5  Rr6  �r7  �r8  hK%�r9  hK%K�r:  �r;  hK�r<  hKhhC   r=  �r>  Rr?  �r@  �rA  hK�rB  hKK�rC  �rD  hK�rE  hKK�rF  �rG  hK�rH  hKK�rI  �rJ  hK�rK  hKhhC   rL  �rM  RrN  �rO  �rP  hK%�rQ  hK%K�rR  �rS  hK�rT  hKhhC   rU  �rV  RrW  �rX  �rY  hK�rZ  hKhhC   r[  �r\  Rr]  �r^  �r_  hK�r`  hKK�ra  �rb  hK�rc  hKK�rd  �re  hK�rf  hKhhC   rg  �rh  Rri  �rj  �rk  hK%�rl  hK%K�rm  �rn  hK�ro  hKhhC   rp  �rq  Rrr  �rs  �rt  hK%�ru  hK%K�rv  �rw  hK�rx  hKhhC   ry  �rz  Rr{  �r|  �r}  hK�r~  hKK�r  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r   �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK%�r  hK%K�r	  �r
  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK%�r   hK%K�r!  �r"  hK�r#  hKK�r$  �r%  hK�r&  hKhhC   r'  �r(  Rr)  �r*  �r+  hK�r,  hKK�r-  �r.  hK�r/  hKhhC   r0  �r1  Rr2  �r3  �r4  hK�r5  hKhhC   r6  �r7  Rr8  �r9  �r:  hK�r;  hKK�r<  �r=  hK%�r>  hK%K�r?  �r@  hK%�rA  hK%K�rB  �rC  hK�rD  hKK�rE  �rF  hK�rG  hKK�rH  �rI  hK�rJ  hKhhC   rK  �rL  RrM  �rN  �rO  hK�rP  hKhhC   rQ  �rR  RrS  �rT  �rU  hK%�rV  hK%K�rW  �rX  hK�rY  hKK�rZ  �r[  hK�r\  hKK�r]  �r^  hK�r_  hKhhC   r`  �ra  Rrb  �rc  �rd  hK�re  hKhhC   rf  �rg  Rrh  �ri  �rj  hK�rk  hKhhC   rl  �rm  Rrn  �ro  �rp  hK�rq  hKK�rr  �rs  hK�rt  hKK�ru  �rv  hK�rw  hKhhC   rx  �ry  Rrz  �r{  �r|  hK%�r}  hK%K�r~  �r  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r   Rr  �r  �r  hK�r  hKK�r  �r  hK%�r  hK%K�r  �r	  hK�r
  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r   �r!  hK�r"  hKK�r#  �r$  hK%�r%  hK%K�r&  �r'  hK�r(  hKK�r)  �r*  hK�r+  hKK�r,  �r-  hK�r.  hKhhC   r/  �r0  Rr1  �r2  �r3  hK�r4  hKhhC   r5  �r6  Rr7  �r8  �r9  hK%�r:  hK%K�r;  �r<  hK%�r=  hK%K�r>  �r?  hK�r@  hKhhC   rA  �rB  RrC  �rD  �rE  hK�rF  hKK�rG  �rH  hK�rI  hKK�rJ  �rK  hK�rL  hKhhC   rM  �rN  RrO  �rP  �rQ  hK�rR  hKhhC   rS  �rT  RrU  �rV  �rW  hK�rX  hKK�rY  �rZ  hK�r[  hKK�r\  �r]  hK%�r^  hK%K�r_  �r`  hK�ra  hKhhC   rb  �rc  Rrd  �re  �rf  hK�rg  hKK�rh  �ri  hK�rj  hKhhC   rk  �rl  Rrm  �rn  �ro  hK�rp  hKK�rq  �rr  hK�rs  hKhhC   rt  �ru  Rrv  �rw  �rx  hK%�ry  hK%K�rz  �r{  hK�r|  hKK�r}  �r~  hK�r  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r   hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r	  hKK�r
  �r  hK%�r  hK%K�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK%�r  hK%K�r  �r   hK�r!  hKK�r"  �r#  hK%�r$  hK%K�r%  �r&  hK�r'  hKhhC   r(  �r)  Rr*  �r+  �r,  hK�r-  hKhhC   r.  �r/  Rr0  �r1  �r2  hK�r3  hKK�r4  �r5  hK�r6  hKK�r7  �r8  hK�r9  hKhhC   r:  �r;  Rr<  �r=  �r>  hK%�r?  hK%K�r@  �rA  hK�rB  hKK�rC  �rD  hK�rE  hKhhC   rF  �rG  RrH  �rI  �rJ  hK�rK  hKK�rL  �rM  hK�rN  hKK�rO  �rP  hK�rQ  hKhhC   rR  �rS  RrT  �rU  �rV  hK�rW  hKhhC   rX  �rY  RrZ  �r[  �r\  hK�r]  hKK�r^  �r_  hK%�r`  hK%K�ra  �rb  hK�rc  hKK�rd  �re  hK�rf  hKhhC   rg  �rh  Rri  �rj  �rk  hK�rl  hKhhC   rm  �rn  Rro  �rp  �rq  hK%�rr  hK%K�rs  �rt  hK�ru  hKK�rv  �rw  hK�rx  hKhhC   ry  �rz  Rr{  �r|  �r}  hK%�r~  hK%K�r  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r   �r  Rr  �r  �r  hK�r  hKhhC   r  �r  Rr  �r	  �r
  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK%�r  hK%K�r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r   hKhhC   r!  �r"  Rr#  �r$  �r%  hK%�r&  hK%K�r'  �r(  hK�r)  hKhhC   r*  �r+  Rr,  �r-  �r.  hK�r/  hKK�r0  �r1  hK�r2  hKK�r3  �r4  hK�r5  hKK�r6  �r7  hK%�r8  hK%K�r9  �r:  hK�r;  hKK�r<  �r=  hK�r>  hKhhC   r?  �r@  RrA  �rB  �rC  hK�rD  hKhhC   rE  �rF  RrG  �rH  �rI  hK�rJ  hKhhC   rK  �rL  RrM  �rN  �rO  hK%�rP  hK%K�rQ  �rR  hK�rS  hKK�rT  �rU  hK�rV  hKK�rW  �rX  hK�rY  hKhhC   rZ  �r[  Rr\  �r]  �r^  hK%�r_  hK%K�r`  �ra  hK�rb  hKK�rc  �rd  hK�re  hKhhC   rf  �rg  Rrh  �ri  �rj  hK�rk  hKK�rl  �rm  hK�rn  hKhhC   ro  �rp  Rrq  �rr  �rs  hK%�rt  hK%K�ru  �rv  hK�rw  hKhhC   rx  �ry  Rrz  �r{  �r|  hK�r}  hKhhC   r~  �r  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r   hK�r  hKK�r  �r  hK�r  hKK�r  �r  hK�r  hKK�r  �r	  hK�r
  hKhhC   r  �r  Rr  �r  �r  hK%�r  hK%K�r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKhhC   r  �r  Rr  �r   �r!  hK�r"  hKK�r#  �r$  hK�r%  hKK�r&  �r'  hK�r(  hKhhC   r)  �r*  Rr+  �r,  �r-  hK%�r.  hK%K�r/  �r0  hK�r1  hKK�r2  �r3  hK�r4  hKK�r5  �r6  hK�r7  hKhhC   r8  �r9  Rr:  �r;  �r<  hK�r=  hKhhC   r>  �r?  Rr@  �rA  �rB  hK%�rC  hK%K�rD  �rE  hK%�rF  hK%K�rG  �rH  hK�rI  hKhhC   rJ  �rK  RrL  �rM  �rN  hK�rO  hKK�rP  �rQ  hK�rR  hKhhC   rS  �rT  RrU  �rV  �rW  hK�rX  hKK�rY  �rZ  hK�r[  hKhhC   r\  �r]  Rr^  �r_  �r`  hK%�ra  hK%K�rb  �rc  hK�rd  hKK�re  �rf  hK�rg  hKhhC   rh  �ri  Rrj  �rk  �rl  hK�rm  hKK�rn  �ro  hK%�rp  hK%K�rq  �rr  hK�rs  hKhhC   rt  �ru  Rrv  �rw  �rx  hK�ry  hKK�rz  �r{  hK�r|  hKK�r}  �r~  hK�r  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r   hK%K�r  �r  hK%�r  hK%K�r  �r  hK�r  hKK�r  �r  hK�r	  hKhhC   r
  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK�r  hKK�r  �r  hK%�r  hK%K�r  �r   hK�r!  hKhhC   r"  �r#  Rr$  �r%  �r&  hK�r'  hKhhC   r(  �r)  Rr*  �r+  �r,  hK�r-  hKhhC   r.  �r/  Rr0  �r1  �r2  hK�r3  hKK�r4  �r5  hK�r6  hKK�r7  �r8  hK�r9  hKhhC   r:  �r;  Rr<  �r=  �r>  hK%�r?  hK%K�r@  �rA  hK%�rB  hK%K�rC  �rD  hK�rE  hKK�rF  �rG  hK�rH  hKhhC   rI  �rJ  RrK  �rL  �rM  hK�rN  hKhhC   rO  �rP  RrQ  �rR  �rS  hK�rT  hKK�rU  �rV  hK�rW  hKK�rX  �rY  hK%�rZ  hK%K�r[  �r\  hK�r]  hKhhC   r^  �r_  Rr`  �ra  �rb  hK�rc  hKK�rd  �re  hK�rf  hKhhC   rg  �rh  Rri  �rj  �rk  hK�rl  hKK�rm  �rn  hK�ro  hKhhC   rp  �rq  Rrr  �rs  �rt  hK�ru  hKK�rv  �rw  hK%�rx  hK%K�ry  �rz  hK�r{  hKhhC   r|  �r}  Rr~  �r  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r   �r  hK�r  hKK�r  �r  hK%�r  hK%K�r  �r  hK�r  hKhhC   r	  �r
  Rr  �r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK%�r  hK%K�r  �r  hK�r  hKhhC   r  �r  Rr   �r!  �r"  hK�r#  hKK�r$  �r%  hK�r&  hKK�r'  �r(  hK�r)  hKhhC   r*  �r+  Rr,  �r-  �r.  hK%�r/  hK%K�r0  �r1  hK�r2  hKhhC   r3  �r4  Rr5  �r6  �r7  hK�r8  hKK�r9  �r:  hK�r;  hKK�r<  �r=  hK�r>  hKhhC   r?  �r@  RrA  �rB  �rC  hK�rD  hKhhC   rE  �rF  RrG  �rH  �rI  hK%�rJ  hK%K�rK  �rL  hK�rM  hKK�rN  �rO  hK�rP  hKK�rQ  �rR  hK�rS  hKK�rT  �rU  hK�rV  hKhhC   rW  �rX  RrY  �rZ  �r[  hK%�r\  hK%K�r]  �r^  hK�r_  hKK�r`  �ra  hK�rb  hKhhC   rc  �rd  Rre  �rf  �rg  hK�rh  hKK�ri  �rj  hK�rk  hKK�rl  �rm  hK�rn  hKhhC   ro  �rp  Rrq  �rr  �rs  hK%�rt  hK%K�ru  �rv  hK�rw  hKhhC   rx  �ry  Rrz  �r{  �r|  hK�r}  hKK�r~  �r  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r 	  hK�r	  hKK�r	  �r	  hK�r	  hKhhC   r	  �r	  Rr	  �r	  �r		  hK�r
	  hKhhC   r	  �r	  Rr	  �r	  �r	  hK�r	  hKK�r	  �r	  hK�r	  hKhhC   r	  �r	  Rr	  �r	  �r	  hK�r	  hKK�r	  �r	  hK�r	  hKhhC   r	  �r	  Rr	  �r 	  �r!	  hK%�r"	  hK%K�r#	  �r$	  hK%�r%	  hK%K�r&	  �r'	  hK�r(	  hKK�r)	  �r*	  hK�r+	  hKK�r,	  �r-	  hK�r.	  hKhhC   r/	  �r0	  Rr1	  �r2	  �r3	  hK�r4	  hKhhC   r5	  �r6	  Rr7	  �r8	  �r9	  hK�r:	  hKK�r;	  �r<	  hK�r=	  hKK�r>	  �r?	  hK�r@	  hKhhC   rA	  �rB	  RrC	  �rD	  �rE	  hK%�rF	  hK%K�rG	  �rH	  hK�rI	  hKhhC   rJ	  �rK	  RrL	  �rM	  �rN	  hK�rO	  hKhhC   rP	  �rQ	  RrR	  �rS	  �rT	  hK�rU	  hKhhC   rV	  �rW	  RrX	  �rY	  �rZ	  hK�r[	  hKK�r\	  �r]	  hK�r^	  hKK�r_	  �r`	  hK%�ra	  hK%K�rb	  �rc	  hK�rd	  hKK�re	  �rf	  hK�rg	  hKhhC   rh	  �ri	  Rrj	  �rk	  �rl	  hK%�rm	  hK%K�rn	  �ro	  hK�rp	  hKhhC   rq	  �rr	  Rrs	  �rt	  �ru	  hK�rv	  hKK�rw	  �rx	  hK�ry	  hKhhC   rz	  �r{	  Rr|	  �r}	  �r~	  hK�r	  hKK�r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK%�r�	  hK%K�r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK%�r�	  hK%K�r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK%�r�	  hK%K�r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK%�r�	  hK%K�r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK%�r�	  hK%K�r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK%�r�	  hK%K�r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK�r�	  hKhhC   r�	  �r�	  Rr�	  �r�	  �r�	  hK�r�	  hKK�r�	  �r�	  hK%�r 
  hK%K�r
  �r
  hK�r
  hKhhC   r
  �r
  Rr
  �r
  �r
  hK�r	
  hKK�r

  �r
  hK�r
  hKhhC   r
  �r
  Rr
  �r
  �r
  hK�r
  hKK�r
  �r
  hK%�r
  hK%K�r
  �r
  hK�r
  hKK�r
  �r
  hK�r
  hKhhC   r
  �r
  Rr
  �r
  �r 
  hK�r!
  hKhhC   r"
  �r#
  Rr$
  �r%
  �r&
  hK�r'
  hKK�r(
  �r)
  hK%�r*
  hK%K�r+
  �r,
  hK�r-
  hKK�r.
  �r/
  hK�r0
  hKhhC   r1
  �r2
  Rr3
  �r4
  �r5
  hK�r6
  hKK�r7
  �r8
  hK�r9
  hKK�r:
  �r;
  hK�r<
  hKhhC   r=
  �r>
  Rr?
  �r@
  �rA
  hK�rB
  hKhhC   rC
  �rD
  RrE
  �rF
  �rG
  hK%�rH
  hK%K�rI
  �rJ
  hK�rK
  hKK�rL
  �rM
  hK�rN
  hKhhC   rO
  �rP
  RrQ
  �rR
  �rS
  hK�rT
  hKK�rU
  �rV
  hK�rW
  hKhhC   rX
  �rY
  RrZ
  �r[
  �r\
  hK%�r]
  hK%K�r^
  �r_
  hK�r`
  hKhhC   ra
  �rb
  Rrc
  �rd
  �re
  hK�rf
  hKK�rg
  �rh
  hK%�ri
  hK%K�rj
  �rk
  hK�rl
  hKhhC   rm
  �rn
  Rro
  �rp
  �rq
  hK�rr
  hKK�rs
  �rt
  hK�ru
  hKhhC   rv
  �rw
  Rrx
  �ry
  �rz
  hK�r{
  hKK�r|
  �r}
  hK�r~
  hKK�r
  �r�
  hK%�r�
  hK%K�r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK�r�
  hKK�r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK�r�
  hKK�r�
  �r�
  hK%�r�
  hK%K�r�
  �r�
  hK%�r�
  hK%K�r�
  �r�
  hK�r�
  hKK�r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK�r�
  hKK�r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK�r�
  hKK�r�
  �r�
  hK%�r�
  hK%K�r�
  �r�
  hK�r�
  hKK�r�
  �r�
  hK�r�
  hKK�r�
  �r�
  hK�r�
  hKK�r�
  �r�
  hK%�r�
  hK%K�r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK�r�
  hKK�r�
  �r�
  hK�r�
  hKK�r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK%�r�
  hK%K�r�
  �r�
  hK�r�
  hKK�r�
  �r�
  hK�r�
  hKhhC   r�
  �r�
  Rr�
  �r�
  �r�
  hK%�r�
  hK%K�r�
  �r�
  hK�r�
  hKK�r   �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK%�r  hK%K�r	  �r
  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKhhC   r  �r  Rr   �r!  �r"  hK�r#  hKK�r$  �r%  hK�r&  hKK�r'  �r(  hK%�r)  hK%K�r*  �r+  hK�r,  hKhhC   r-  �r.  Rr/  �r0  �r1  hK�r2  hKK�r3  �r4  hK�r5  hKhhC   r6  �r7  Rr8  �r9  �r:  hK�r;  hKK�r<  �r=  hK�r>  hKhhC   r?  �r@  RrA  �rB  �rC  hK%�rD  hK%K�rE  �rF  hK�rG  hKhhC   rH  �rI  RrJ  �rK  �rL  hK�rM  hKK�rN  �rO  hK�rP  hKhhC   rQ  �rR  RrS  �rT  �rU  hK�rV  hKK�rW  �rX  hK%�rY  hK%K�rZ  �r[  hK�r\  hKhhC   r]  �r^  Rr_  �r`  �ra  hK�rb  hKK�rc  �rd  hK�re  hKK�rf  �rg  hK�rh  hKhhC   ri  �rj  Rrk  �rl  �rm  hK%�rn  hK%K�ro  �rp  hK�rq  hKK�rr  �rs  hK�rt  hKhhC   ru  �rv  Rrw  �rx  �ry  hK%�rz  hK%K�r{  �r|  hK�r}  hKhhC   r~  �r  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r   hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r	  hK�r
  hKK�r  �r  hK�r  hKK�r  �r  hK%�r  hK%K�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK%�r  hK%K�r  �r  hK�r  hKK�r   �r!  hK�r"  hKhhC   r#  �r$  Rr%  �r&  �r'  hK�r(  hKhhC   r)  �r*  Rr+  �r,  �r-  hK�r.  hKhhC   r/  �r0  Rr1  �r2  �r3  hK�r4  hKhhC   r5  �r6  Rr7  �r8  �r9  hK�r:  hKK�r;  �r<  hK�r=  hKK�r>  �r?  hK%�r@  hK%K�rA  �rB  hK�rC  hKhhC   rD  �rE  RrF  �rG  �rH  hK%�rI  hK%K�rJ  �rK  hK�rL  hKK�rM  �rN  hK�rO  hKK�rP  �rQ  hK�rR  hKhhC   rS  �rT  RrU  �rV  �rW  hK�rX  hKK�rY  �rZ  hK�r[  hKhhC   r\  �r]  Rr^  �r_  �r`  hK�ra  hKhhC   rb  �rc  Rrd  �re  �rf  hK%�rg  hK%K�rh  �ri  hK�rj  hKK�rk  �rl  hK�rm  hKK�rn  �ro  hK�rp  hKK�rq  �rr  hK�rs  hKhhC   rt  �ru  Rrv  �rw  �rx  hK%�ry  hK%K�rz  �r{  hK�r|  hKhhC   r}  �r~  Rr  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r   hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK�r	  hKK�r
  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK%�r  hK%K�r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK%�r  hK%K�r  �r   hK�r!  hKK�r"  �r#  hK�r$  hKhhC   r%  �r&  Rr'  �r(  �r)  hK%�r*  hK%K�r+  �r,  hK�r-  hKhhC   r.  �r/  Rr0  �r1  �r2  hK�r3  hKK�r4  �r5  hK�r6  hKhhC   r7  �r8  Rr9  �r:  �r;  hK�r<  hKK�r=  �r>  hK�r?  hKhhC   r@  �rA  RrB  �rC  �rD  hK�rE  hKK�rF  �rG  hK%�rH  hK%K�rI  �rJ  hK�rK  hKK�rL  �rM  hK�rN  hKhhC   rO  �rP  RrQ  �rR  �rS  hK%�rT  hK%K�rU  �rV  hK�rW  hKhhC   rX  �rY  RrZ  �r[  �r\  hK�r]  hKK�r^  �r_  hK�r`  hKhhC   ra  �rb  Rrc  �rd  �re  hK�rf  hKK�rg  �rh  hK�ri  hKK�rj  �rk  hK�rl  hKhhC   rm  �rn  Rro  �rp  �rq  hK�rr  hKhhC   rs  �rt  Rru  �rv  �rw  hK�rx  hKK�ry  �rz  hK%�r{  hK%K�r|  �r}  hK%�r~  hK%K�r  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r   �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r	  �r
  hK�r  hKK�r  �r  hK%�r  hK%K�r  �r  hK�r  hKK�r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKhhC   r  �r  Rr   �r!  �r"  hK%�r#  hK%K�r$  �r%  hK�r&  hKhhC   r'  �r(  Rr)  �r*  �r+  hK�r,  hKK�r-  �r.  hK�r/  hKK�r0  �r1  hK�r2  hKhhC   r3  �r4  Rr5  �r6  �r7  hK%�r8  hK%K�r9  �r:  hK%�r;  hK%K�r<  �r=  hK�r>  hKhhC   r?  �r@  RrA  �rB  �rC  hK�rD  hKK�rE  �rF  hK�rG  hKhhC   rH  �rI  RrJ  �rK  �rL  hK�rM  hKK�rN  �rO  hK%�rP  hK%K�rQ  �rR  hK�rS  hKK�rT  �rU  hK�rV  hKK�rW  �rX  hK�rY  hKhhC   rZ  �r[  Rr\  �r]  �r^  hK�r_  hKhhC   r`  �ra  Rrb  �rc  �rd  hK%�re  hK%K�rf  �rg  hK�rh  hKK�ri  �rj  hK�rk  hKhhC   rl  �rm  Rrn  �ro  �rp  hK�rq  hKK�rr  �rs  hK�rt  hKhhC   ru  �rv  Rrw  �rx  �ry  hK�rz  hKK�r{  �r|  hK�r}  hKhhC   r~  �r  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r   hK%�r  hK%K�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r	  hK�r
  hKK�r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK%�r  hK%K�r   �r!  hK�r"  hKK�r#  �r$  hK�r%  hKhhC   r&  �r'  Rr(  �r)  �r*  hK%�r+  hK%K�r,  �r-  hK�r.  hKK�r/  �r0  hK�r1  hKhhC   r2  �r3  Rr4  �r5  �r6  hK�r7  hKK�r8  �r9  hK%�r:  hK%K�r;  �r<  hK�r=  hKK�r>  �r?  hK�r@  hKhhC   rA  �rB  RrC  �rD  �rE  hK�rF  hKhhC   rG  �rH  RrI  �rJ  �rK  hK�rL  hKhhC   rM  �rN  RrO  �rP  �rQ  hK�rR  hKK�rS  �rT  hK�rU  hKhhC   rV  �rW  RrX  �rY  �rZ  hK�r[  hKK�r\  �r]  hK%�r^  hK%K�r_  �r`  hK�ra  hKK�rb  �rc  hK%�rd  hK%K�re  �rf  hK�rg  hKK�rh  �ri  hK�rj  hKhhC   rk  �rl  Rrm  �rn  �ro  hK�rp  hKhhC   rq  �rr  Rrs  �rt  �ru  hK�rv  hKK�rw  �rx  hK�ry  hKK�rz  �r{  hK%�r|  hK%K�r}  �r~  hK�r  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr   �r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r	  hKK�r
  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK%�r  hK%K�r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK%�r  hK%K�r  �r   hK�r!  hKhhC   r"  �r#  Rr$  �r%  �r&  hK�r'  hKK�r(  �r)  hK�r*  hKK�r+  �r,  hK�r-  hKhhC   r.  �r/  Rr0  �r1  �r2  hK�r3  hKhhC   r4  �r5  Rr6  �r7  �r8  hK�r9  hKK�r:  �r;  hK�r<  hKhhC   r=  �r>  Rr?  �r@  �rA  hK�rB  hKK�rC  �rD  hK%�rE  hK%K�rF  �rG  hK%�rH  hK%K�rI  �rJ  hK�rK  hKhhC   rL  �rM  RrN  �rO  �rP  hK�rQ  hKK�rR  �rS  hK�rT  hKhhC   rU  �rV  RrW  �rX  �rY  hK�rZ  hKK�r[  �r\  hK�r]  hKhhC   r^  �r_  Rr`  �ra  �rb  hK�rc  hKK�rd  �re  hK%�rf  hK%K�rg  �rh  hK�ri  hKhhC   rj  �rk  Rrl  �rm  �rn  hK�ro  hKK�rp  �rq  e(hK�rr  hKhhC   rs  �rt  Rru  �rv  �rw  hK�rx  hKK�ry  �rz  hK�r{  hKK�r|  �r}  hK%�r~  hK%K�r  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r   �r  hK%�r  hK%K�r  �r  hK�r  hKhhC   r  �r  Rr  �r	  �r
  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK�r  hKK�r  �r  hK%�r  hK%K�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK%�r   hK%K�r!  �r"  hK�r#  hKK�r$  �r%  hK�r&  hKK�r'  �r(  hK�r)  hKhhC   r*  �r+  Rr,  �r-  �r.  hK�r/  hKK�r0  �r1  hK%�r2  hK%K�r3  �r4  hK�r5  hKhhC   r6  �r7  Rr8  �r9  �r:  hK�r;  hKhhC   r<  �r=  Rr>  �r?  �r@  hK�rA  hKK�rB  �rC  hK�rD  hKhhC   rE  �rF  RrG  �rH  �rI  hK%�rJ  hK%K�rK  �rL  hK�rM  hKhhC   rN  �rO  RrP  �rQ  �rR  hK�rS  hKK�rT  �rU  hK�rV  hKK�rW  �rX  hK%�rY  hK%K�rZ  �r[  hK�r\  hKhhC   r]  �r^  Rr_  �r`  �ra  hK�rb  hKK�rc  �rd  hK�re  hKhhC   rf  �rg  Rrh  �ri  �rj  hK�rk  hKK�rl  �rm  hK�rn  hKK�ro  �rp  hK�rq  hKK�rr  �rs  hK�rt  hKhhC   ru  �rv  Rrw  �rx  �ry  hK�rz  hKhhC   r{  �r|  Rr}  �r~  �r  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r   hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r	  hK�r
  hKK�r  �r  hK%�r  hK%K�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r   �r!  Rr"  �r#  �r$  hK�r%  hKK�r&  �r'  hK%�r(  hK%K�r)  �r*  hK�r+  hKK�r,  �r-  hK%�r.  hK%K�r/  �r0  hK�r1  hKK�r2  �r3  hK�r4  hKhhC   r5  �r6  Rr7  �r8  �r9  hK�r:  hKhhC   r;  �r<  Rr=  �r>  �r?  hK�r@  hKK�rA  �rB  hK%�rC  hK%K�rD  �rE  hK�rF  hKK�rG  �rH  hK�rI  hKhhC   rJ  �rK  RrL  �rM  �rN  hK�rO  hKhhC   rP  �rQ  RrR  �rS  �rT  hK�rU  hKK�rV  �rW  hK�rX  hKhhC   rY  �rZ  Rr[  �r\  �r]  hK�r^  hKK�r_  �r`  hK%�ra  hK%K�rb  �rc  hK�rd  hKhhC   re  �rf  Rrg  �rh  �ri  hK�rj  hKK�rk  �rl  hK�rm  hKK�rn  �ro  hK�rp  hKhhC   rq  �rr  Rrs  �rt  �ru  hK%�rv  hK%K�rw  �rx  hK�ry  hKhhC   rz  �r{  Rr|  �r}  �r~  hK�r  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r   hKhhC   r  �r  Rr  �r  �r  hK�r  hKK�r  �r  hK�r	  hKhhC   r
  �r  Rr  �r  �r  hK%�r  hK%K�r  �r  hK�r  hKK�r  �r  hK%�r  hK%K�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKhhC   r  �r   Rr!  �r"  �r#  hK�r$  hKK�r%  �r&  hK�r'  hKK�r(  �r)  hK�r*  hKK�r+  �r,  hK%�r-  hK%K�r.  �r/  hK�r0  hKhhC   r1  �r2  Rr3  �r4  �r5  hK�r6  hKhhC   r7  �r8  Rr9  �r:  �r;  hK�r<  hKhhC   r=  �r>  Rr?  �r@  �rA  hK%�rB  hK%K�rC  �rD  hK�rE  hKK�rF  �rG  hK�rH  hKK�rI  �rJ  hK�rK  hKhhC   rL  �rM  RrN  �rO  �rP  hK�rQ  hKhhC   rR  �rS  RrT  �rU  �rV  hK%�rW  hK%K�rX  �rY  hK�rZ  hKhhC   r[  �r\  Rr]  �r^  �r_  hK�r`  hKK�ra  �rb  hK�rc  hKK�rd  �re  hK�rf  hKK�rg  �rh  hK�ri  hKK�rj  �rk  hK�rl  hKhhC   rm  �rn  Rro  �rp  �rq  hK%�rr  hK%K�rs  �rt  hK�ru  hKhhC   rv  �rw  Rrx  �ry  �rz  hK�r{  hKK�r|  �r}  hK�r~  hKhhC   r  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK%�r�  hK%K�r   �r  hK�r  hKK�r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r	  �r
  Rr  �r  �r  hK%�r  hK%K�r  �r  hK�r  hKK�r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r  hKhhC   r  �r  Rr  �r  �r  hK�r   hKK�r!  �r"  hK�r#  hKK�r$  �r%  hK�r&  hKK�r'  �r(  hK%�r)  hK%K�r*  �r+  hK�r,  hKhhC   r-  �r.  Rr/  �r0  �r1  hK�r2  hKhhC   r3  �r4  Rr5  �r6  �r7  hK�r8  hKK�r9  �r:  hK�r;  hKK�r<  �r=  hK�r>  hKhhC   r?  �r@  RrA  �rB  �rC  hK%�rD  hK%K�rE  �rF  hK�rG  hKhhC   rH  �rI  RrJ  �rK  �rL  hK�rM  hKhhC   rN  �rO  RrP  �rQ  �rR  hK�rS  hKK�rT  �rU  hK�rV  hKhhC   rW  �rX  RrY  �rZ  �r[  hK%�r\  hK%K�r]  �r^  hK�r_  hKK�r`  �ra  hK�rb  hKhhC   rc  �rd  Rre  �rf  �rg  hK�rh  hKK�ri  �rj  hK�rk  hKK�rl  �rm  hK%�rn  hK%K�ro  �rp  hK�rq  hKhhC   rr  �rs  Rrt  �ru  �rv  hK�rw  hKhhC   rx  �ry  Rrz  �r{  �r|  hK%�r}  hK%K�r~  �r  hK�r�  hKK�r�  �r�  hK�r�  hKhhC   r�  �r�  Rr�  �r�  �r�  hK�r�  hKK�r�  �r�  e.