�]q (]q(]q(X   Normsq]q(X   Oblq]q(X   Movedq]q(X   Colourq	X   rq
e]q(X   ShapeqX   circleqe]q(X   ZoneqX   3qe]q(X   Movedq]q(h	X   bqe]q(hX   squareqe]q(hX   1qe]q(X	   Next-Moveq]q(h	he]q(hX   triangleqeeee]q(hX   2qee]q (X   Perq!]q"(X   Actionq#X   putdownq$e]q%(h	h
e]q&(hX   triangleq'e]q((X   PerZoneq)heee]q*(h]q+(h]q,(h]q-(h	h
e]q.(hhe]q/(hhe]q0(h]q1(h	he]q2(hhe]q3(hhe]q4(h]q5(h	he]q6(hheeee]q7(hhee]q8(h!]q9(h#h$e]q:(h	he]q;(hX   circleq<e]q=(h)heeeh*h*]q>(h]q?(h]q@(h]qA(h	h
e]qB(hhe]qC(hhe]qD(h]qE(h	he]qF(hhe]qG(hhe]qH(h]qI(h	he]qJ(hheeee]qK(hhee]qL(h!]qM(h#h$e]qN(h	he]qO(hh<e]qP(h)heeeh>h>]qQ(h]qR(h]qS(h]qT(h	h
e]qU(hhe]qV(hhe]qW(h]qX(h	he]qY(hhe]qZ(hhe]q[(h]q\(h	he]q](hheeee]q^(hhee]q_(h!]q`(h#h$e]qa(h	he]qb(hh<e]qc(h)heee]qd(h]qe(h]qf(h]qg(h	h
e]qh(hhe]qi(hhe]qj(h]qk(h	he]ql(hhe]qm(hhe]qn(h]qo(h	he]qp(hheeee]qq(hhee]qr(h!]qs(h#h$e]qt(h	he]qu(hh<e]qv(h)heeehdhdhdhdhdhd]qw(h]qx(h]qy(h]qz(h	h
e]q{(hhe]q|(hhe]q}(h]q~(h	he]q(hhe]q�(hhe]q�(h]q�(h	he]q�(hheeee]q�(hhee]q�(h!]q�(h#h$e]q�(h	X   anyq�e]q�(hX   squareq�e]q�(h)heee]q�(h]q�(h]q�(h]q�(h	h
e]q�(hhe]q�(hhe]q�(h]q�(h	he]q�(hhe]q�(hhe]q�(h]q�(h	he]q�(hheeee]q�(hhee]q�(h!]q�(h#h$e]q�(h	h�e]q�(hh�e]q�(h)heee]q�(h]q�(h]q�(h]q�(h	h
e]q�(hhe]q�(hhe]q�(h]q�(h	he]q�(hhe]q�(hhe]q�(h]q�(h	he]q�(hheeee]q�(hhee]q�(h!]q�(h#h$e]q�(h	h�e]q�(hh�e]q�(h)heeeh�h�]q�(h]q�(h]q�(h]q�(h	h
e]q�(hhe]q�(hhe]q�(h]q�(h	he]q�(hhe]q�(hhe]q�(h]q�(h	he]q�(hheeee]q�(hhee]q�(h!]q�(h#h$e]q�(h	h�e]q�(hh�e]q�(h)heee]q�(h]q�(h]q�(h]q�(h	h
e]q�(hhe]q�(hhe]q�(h]q�(h	he]q�(hh�e]q�(hhe]q�(h]q�(h	he]q�(hheeee]q�(hhee]q�(h!]q�(h#h$e]q�(h	h�e]q�(hh�e]q�(h)heee]q�(h]q�(h]q�(h]q�(h	h
e]q�(hhe]q�(hhe]q�(h]q�(h	he]q�(hh�e]q�(hhe]q�(h]q�(h	he]q�(hheeee]q�(hhee]q�(h!]q�(h#h$e]q�(h	h�e]q�(hh�e]q�(h)heee]q�(h]q�(h]q�(h]q�(h	h
e]q�(hhe]q�(hhe]q�(h]q�(h	he]q�(hh�e]q�(hhe]q�(h]q�(h	he]q�(hX   triangleq�eeee]q�(hhee]q�(h!]q�(h#h$e]q�(h	h�e]q�(hh�e]q�(h)heeeh�h�h�]q�(h]r   (h]r  (h]r  (h	h
e]r  (hhe]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r	  (h]r
  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	h�e]r  (hh�e]r  (h)heee]r  (h]r  (h]r  (h]r  (h	h
e]r  (hhe]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�eeee]r  (hhee]r   (h!]r!  (h#h$e]r"  (h	h�e]r#  (hh�e]r$  (h)heee]r%  (h]r&  (h]r'  (h]r(  (h	h
e]r)  (hhe]r*  (hhe]r+  (h]r,  (h	he]r-  (hh�e]r.  (hhe]r/  (h]r0  (h	he]r1  (hh�eeee]r2  (hhee]r3  (h!]r4  (h#h$e]r5  (h	h�e]r6  (hh�e]r7  (h)heeej%  ]r8  (h]r9  (h]r:  (h]r;  (h	h
e]r<  (hhe]r=  (hhe]r>  (h]r?  (h	he]r@  (hh�e]rA  (hhe]rB  (h]rC  (h	he]rD  (hh�eeee]rE  (hhee]rF  (h!]rG  (h#h$e]rH  (h	h�e]rI  (hh�e]rJ  (h)heeej8  j8  j8  ]rK  (h]rL  (h]rM  (h]rN  (h	h
e]rO  (hhe]rP  (hhe]rQ  (h]rR  (h	he]rS  (hh�e]rT  (hhe]rU  (h]rV  (h	he]rW  (hh�eeee]rX  (hhee]rY  (h!]rZ  (h#h$e]r[  (h	h�e]r\  (hh�e]r]  (h)heee]r^  (h]r_  (h]r`  (h]ra  (h	h
e]rb  (hhe]rc  (hhe]rd  (h]re  (h	he]rf  (hh�e]rg  (hhe]rh  (h]ri  (h	he]rj  (hh�eeee]rk  (hhee]rl  (h!]rm  (h#h$e]rn  (h	h�e]ro  (hh�e]rp  (h)heee]rq  (h]rr  (h]rs  (h]rt  (h	h
e]ru  (hhe]rv  (hhe]rw  (h]rx  (h	he]ry  (hh�e]rz  (hhe]r{  (h]r|  (h	he]r}  (hh�eeee]r~  (hhee]r  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejq  jq  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hhe]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hhe]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hhe]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hhe]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hhe]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hhe]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hhe]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r   (h]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	h�e]r  (hh�e]r  (h)heeej�  j�  j�  j�  j�  j�  j�  ]r	  (h]r
  (h]r  (h]r  (h	h
e]r  (hhe]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	h�e]r  (hh�e]r  (h)heee]r  (h]r  (h]r  (h]r  (h	h
e]r   (hhe]r!  (hhe]r"  (h]r#  (h	he]r$  (hh�e]r%  (hhe]r&  (h]r'  (h	he]r(  (hh�eeee]r)  (hhee]r*  (h!]r+  (h#h$e]r,  (h	h�e]r-  (hh�e]r.  (h)heee]r/  (h]r0  (h]r1  (h]r2  (h	h
e]r3  (hhe]r4  (hhe]r5  (h]r6  (h	he]r7  (hh�e]r8  (hhe]r9  (h]r:  (h	he]r;  (hh�eeee]r<  (hhee]r=  (h!]r>  (h#h$e]r?  (h	h�e]r@  (hh�e]rA  (h)heee]rB  (h]rC  (h]rD  (h]rE  (h	h
e]rF  (hhe]rG  (hhe]rH  (h]rI  (h	he]rJ  (hh�e]rK  (hhe]rL  (h]rM  (h	he]rN  (hh�eeee]rO  (hhee]rP  (h!]rQ  (h#h$e]rR  (h	h
e]rS  (hh<e]rT  (h)heee]rU  (h]rV  (h]rW  (h]rX  (h	h
e]rY  (hhe]rZ  (hhe]r[  (h]r\  (h	he]r]  (hh�e]r^  (hhe]r_  (h]r`  (h	he]ra  (hh�eeee]rb  (hhee]rc  (h!]rd  (h#h$e]re  (h	h
e]rf  (hh<e]rg  (h)heee]rh  (h]ri  (h]rj  (h]rk  (h	h
e]rl  (hhe]rm  (hhe]rn  (h]ro  (h	he]rp  (hh�e]rq  (hhe]rr  (h]rs  (h	he]rt  (hh�eeee]ru  (hhee]rv  (h!]rw  (h#h$e]rx  (h	h
e]ry  (hh<e]rz  (h)heeejh  ]r{  (h]r|  (h]r}  (h]r~  (h	h
e]r  (hhe]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh<e]r�  (h)heeej{  j{  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh<e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh<e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eeej�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eeej�  ]r   (h]r  (h]r  (h]r  (h	h
e]r  (hh<e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r	  (hhe]r
  (h]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	h
e]r  (hh�e]r  (h)h�eee]r  (h]r  (h]r  (h]r  (h	h
e]r  (hh<e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�eeee]r   (hhee]r!  (h!]r"  (h#h$e]r#  (h	h
e]r$  (hh<e]r%  (h)h�eeej  j  j  j  ]r&  (h]r'  (h]r(  (h]r)  (h	h
e]r*  (hh<e]r+  (hhe]r,  (h]r-  (h	he]r.  (hh�e]r/  (hhe]r0  (h]r1  (h	h�e]r2  (hh�eeee]r3  (hhee]r4  (h!]r5  (h#h$e]r6  (h	h
e]r7  (hh<e]r8  (h)heee]r9  (h]r:  (h]r;  (h]r<  (h	h
e]r=  (hh<e]r>  (hhe]r?  (h]r@  (h	he]rA  (hh�e]rB  (hhe]rC  (h]rD  (h	h�e]rE  (hh�eeee]rF  (hhee]rG  (h!]rH  (h#h$e]rI  (h	h
e]rJ  (hh<e]rK  (h)heeej9  j9  j9  j9  ]rL  (h]rM  (h]rN  (h]rO  (h	h
e]rP  (hh<e]rQ  (hhe]rR  (h]rS  (h	he]rT  (hh�e]rU  (hhe]rV  (h]rW  (h	h�e]rX  (hh�eeee]rY  (hhee]rZ  (h!]r[  (h#h$e]r\  (h	h�e]r]  (hh�e]r^  (h)h�eee]r_  (h]r`  (h]ra  (h]rb  (h	h
e]rc  (hh<e]rd  (hhe]re  (h]rf  (h	he]rg  (hh�e]rh  (hhe]ri  (h]rj  (h	h�e]rk  (hh�eeee]rl  (hhee]rm  (h!]rn  (h#h$e]ro  (h	h�e]rp  (hh�e]rq  (h)h�eee]rr  (h]rs  (h]rt  (h]ru  (h	h
e]rv  (hh<e]rw  (hhe]rx  (h]ry  (h	he]rz  (hh�e]r{  (hhe]r|  (h]r}  (h	h�e]r~  (hh�eeee]r  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)h�eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)h�eeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r   (hhe]r  (h]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	h
e]r  (hh�e]r	  (h)h�eeej�  j�  j�  ]r
  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	h
e]r  (hh�e]r  (h)h�eee]r  (h]r  (h]r  (h]r   (h	h�e]r!  (hh�e]r"  (hhe]r#  (h]r$  (h	he]r%  (hh�e]r&  (hhe]r'  (h]r(  (h	h�e]r)  (hh�eeee]r*  (hhee]r+  (h!]r,  (h#h$e]r-  (h	h
e]r.  (hh�e]r/  (h)h�eeej  j  ]r0  (h]r1  (h]r2  (h]r3  (h	h�e]r4  (hh�e]r5  (hhe]r6  (h]r7  (h	he]r8  (hh�e]r9  (hhe]r:  (h]r;  (h	h�e]r<  (hh�eeee]r=  (hhee]r>  (h!]r?  (h#h$e]r@  (h	h
e]rA  (hh�e]rB  (h)h�eeej0  ]rC  (h]rD  (h]rE  (h]rF  (h	h�e]rG  (hh�e]rH  (hhe]rI  (h]rJ  (h	he]rK  (hh�e]rL  (hhe]rM  (h]rN  (h	h�e]rO  (hh�eeee]rP  (hhee]rQ  (h!]rR  (h#h$e]rS  (h	h
e]rT  (hh�e]rU  (h)h�eee]rV  (h]rW  (h]rX  (h]rY  (h	h�e]rZ  (hh�e]r[  (hhe]r\  (h]r]  (h	he]r^  (hh�e]r_  (hhe]r`  (h]ra  (h	h�e]rb  (hh�eeee]rc  (hhee]rd  (h!]re  (h#h$e]rf  (h	h
e]rg  (hh�e]rh  (h)h�eee]ri  (h]rj  (h]rk  (h]rl  (h	h�e]rm  (hh�e]rn  (hhe]ro  (h]rp  (h	he]rq  (hh�e]rr  (hhe]rs  (h]rt  (h	h�e]ru  (hh�eeee]rv  (hhee]rw  (h!]rx  (h#h$e]ry  (h	h
e]rz  (hh�e]r{  (h)h�eee]r|  (h]r}  (h]r~  (h]r  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heeej|  j|  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)h�eeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)h�eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r   (h)heeej�  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r	  (hh�e]r
  (hhe]r  (h]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	he]r  (hh<e]r  (h)heee]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r   (hh�eeee]r!  (hhee]r"  (h!]r#  (h#h$e]r$  (h	he]r%  (hh<e]r&  (h)heeej  j  ]r'  (h]r(  (h]r)  (h]r*  (h	h�e]r+  (hh�e]r,  (hhe]r-  (h]r.  (h	he]r/  (hh�e]r0  (hhe]r1  (h]r2  (h	h�e]r3  (hh�eeee]r4  (hhee]r5  (h!]r6  (h#h$e]r7  (h	he]r8  (hh<e]r9  (h)heeej'  ]r:  (h]r;  (h]r<  (h]r=  (h	h�e]r>  (hh�e]r?  (hhe]r@  (h]rA  (h	he]rB  (hh�e]rC  (hhe]rD  (h]rE  (h	h�e]rF  (hh�eeee]rG  (hhee]rH  (h!]rI  (h#h$e]rJ  (h	h
e]rK  (hh<e]rL  (h)heee]rM  (h]rN  (h]rO  (h]rP  (h	h�e]rQ  (hh�e]rR  (hhe]rS  (h]rT  (h	he]rU  (hh�e]rV  (hhe]rW  (h]rX  (h	h�e]rY  (hh�eeee]rZ  (hhee]r[  (h!]r\  (h#h$e]r]  (h	h
e]r^  (hh<e]r_  (h)heeejM  ]r`  (h]ra  (h]rb  (h]rc  (h	h�e]rd  (hh�e]re  (hhe]rf  (h]rg  (h	he]rh  (hh�e]ri  (hhe]rj  (h]rk  (h	h�e]rl  (hh�eeee]rm  (hhee]rn  (h!]ro  (h#h$e]rp  (h	h
e]rq  (hh�e]rr  (h)heee]rs  (h]rt  (h]ru  (h]rv  (h	h�e]rw  (hh�e]rx  (hhe]ry  (h]rz  (h	he]r{  (hh�e]r|  (hhe]r}  (h]r~  (h	h�e]r  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	X   gr�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)h�eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r   (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r	  (h	j�  e]r
  (hh�e]r  (h)heee]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej  j  j  j  j  j  ]r  (h]r   (h]r!  (h]r"  (h	h�e]r#  (hh�e]r$  (hhe]r%  (h]r&  (h	he]r'  (hh�e]r(  (hhe]r)  (h]r*  (h	h�e]r+  (hh�eeee]r,  (hhee]r-  (h!]r.  (h#h$e]r/  (h	j�  e]r0  (hh�e]r1  (h)heeej  j  j  j  ]r2  (h]r3  (h]r4  (h]r5  (h	h�e]r6  (hh�e]r7  (hhe]r8  (h]r9  (h	he]r:  (hh�e]r;  (hhe]r<  (h]r=  (h	h�e]r>  (hh�eeee]r?  (hhee]r@  (h!]rA  (h#h$e]rB  (h	j�  e]rC  (hh�e]rD  (h)heeej2  j2  ]rE  (h]rF  (h]rG  (h]rH  (h	h�e]rI  (hh�e]rJ  (hhe]rK  (h]rL  (h	he]rM  (hh�e]rN  (hhe]rO  (h]rP  (h	he]rQ  (hh�eeee]rR  (hhee]rS  (h!]rT  (h#h$e]rU  (h	j�  e]rV  (hh�e]rW  (h)heeejE  ]rX  (h]rY  (h]rZ  (h]r[  (h	h�e]r\  (hh�e]r]  (hhe]r^  (h]r_  (h	he]r`  (hh�e]ra  (hhe]rb  (h]rc  (h	he]rd  (hh�eeee]re  (hhee]rf  (h!]rg  (h#h$e]rh  (h	j�  e]ri  (hh�e]rj  (h)heee]rk  (h]rl  (h]rm  (h]rn  (h	h�e]ro  (hh�e]rp  (hhe]rq  (h]rr  (h	he]rs  (hh�e]rt  (hhe]ru  (h]rv  (h	he]rw  (hh�eeee]rx  (hhee]ry  (h!]rz  (h#h$e]r{  (h	j�  e]r|  (hh�e]r}  (h)heeejk  ]r~  (h]r  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej~  j~  j~  j~  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r   (h	h
e]r  (hh�e]r  (h)h�eeej�  j�  j�  j�  j�  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r	  (h]r
  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	h
e]r  (hh�e]r  (h)heeej  j  j  j  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r   (h]r!  (h	he]r"  (hh�eeee]r#  (hhee]r$  (h!]r%  (h#h$e]r&  (h	h
e]r'  (hh�e]r(  (h)heeej  j  ]r)  (h]r*  (h]r+  (h]r,  (h	h�e]r-  (hh�e]r.  (hhe]r/  (h]r0  (h	he]r1  (hh�e]r2  (hhe]r3  (h]r4  (h	he]r5  (hh�eeee]r6  (hhee]r7  (h!]r8  (h#h$e]r9  (h	he]r:  (hh�e]r;  (h)heee]r<  (h]r=  (h]r>  (h]r?  (h	h�e]r@  (hh�e]rA  (hhe]rB  (h]rC  (h	he]rD  (hh�e]rE  (hhe]rF  (h]rG  (h	he]rH  (hh�eeee]rI  (hhee]rJ  (h!]rK  (h#h$e]rL  (h	he]rM  (hh�e]rN  (h)heeej<  j<  j<  j<  ]rO  (h]rP  (h]rQ  (h]rR  (h	h�e]rS  (hh�e]rT  (hhe]rU  (h]rV  (h	he]rW  (hh�e]rX  (hhe]rY  (h]rZ  (h	he]r[  (hh�eeee]r\  (hhee]r]  (h!]r^  (h#h$e]r_  (h	he]r`  (hh<e]ra  (h)heee]rb  (h]rc  (h]rd  (h]re  (h	h�e]rf  (hh�e]rg  (hhe]rh  (h]ri  (h	he]rj  (hh�e]rk  (hhe]rl  (h]rm  (h	he]rn  (hh�eeee]ro  (hhee]rp  (h!]rq  (h#h$e]rr  (h	he]rs  (hh<e]rt  (h)heeejb  jb  jb  ]ru  (h]rv  (h]rw  (h]rx  (h	h�e]ry  (hh�e]rz  (hhe]r{  (h]r|  (h	he]r}  (hh�e]r~  (hhe]r  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r   (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r	  (h#h$e]r
  (h	he]r  (hh�e]r  (h)heee]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	he]r  (hh<e]r  (h)heee]r   (h]r!  (h]r"  (h]r#  (h	h�e]r$  (hh<e]r%  (hhe]r&  (h]r'  (h	he]r(  (hh�e]r)  (hhe]r*  (h]r+  (h	he]r,  (hh�eeee]r-  (hhee]r.  (h!]r/  (h#h$e]r0  (h	he]r1  (hh<e]r2  (h)heee]r3  (h]r4  (h]r5  (h]r6  (h	h�e]r7  (hh<e]r8  (hhe]r9  (h]r:  (h	he]r;  (hh�e]r<  (hhe]r=  (h]r>  (h	he]r?  (hh�eeee]r@  (hhee]rA  (h!]rB  (h#h$e]rC  (h	he]rD  (hh<e]rE  (h)heeej3  j3  j3  ]rF  (h]rG  (h]rH  (h]rI  (h	h�e]rJ  (hh�e]rK  (hhe]rL  (h]rM  (h	he]rN  (hh�e]rO  (hhe]rP  (h]rQ  (h	he]rR  (hh�eeee]rS  (hhee]rT  (h!]rU  (h#h$e]rV  (h	he]rW  (hh<e]rX  (h)heee]rY  (h]rZ  (h]r[  (h]r\  (h	h�e]r]  (hh�e]r^  (hhe]r_  (h]r`  (h	he]ra  (hh�e]rb  (hhe]rc  (h]rd  (h	he]re  (hh�eeee]rf  (hhee]rg  (h!]rh  (h#h$e]ri  (h	h�e]rj  (hh�e]rk  (h)heeejY  jY  ]rl  (h]rm  (h]rn  (h]ro  (h	h�e]rp  (hh�e]rq  (hhe]rr  (h]rs  (h	he]rt  (hh�e]ru  (hhe]rv  (h]rw  (h	he]rx  (hh�eeee]ry  (hhee]rz  (h!]r{  (h#h$e]r|  (h	h�e]r}  (hh�e]r~  (h)heee]r  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej  j  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r 	  (h#h$e]r	  (h	h�e]r	  (hh�e]r	  (h)heeej�  j�  ]r	  (h]r	  (h]r	  (h]r	  (h	h�e]r	  (hh<e]r		  (hhe]r
	  (h]r	  (h	he]r	  (hh�e]r	  (hhe]r	  (h]r	  (h	he]r	  (hh�eeee]r	  (hhee]r	  (h!]r	  (h#h$e]r	  (h	h�e]r	  (hh�e]r	  (h)heeej	  ]r	  (h]r	  (h]r	  (h]r	  (h	h�e]r	  (hh<e]r	  (hhe]r	  (h]r	  (h	he]r	  (hh�e]r 	  (hhe]r!	  (h]r"	  (h	he]r#	  (hh�eeee]r$	  (hhee]r%	  (h!]r&	  (h#h$e]r'	  (h	h�e]r(	  (hh�e]r)	  (h)heee]r*	  (h]r+	  (h]r,	  (h]r-	  (h	h�e]r.	  (hh<e]r/	  (hhe]r0	  (h]r1	  (h	he]r2	  (hh�e]r3	  (hhe]r4	  (h]r5	  (h	he]r6	  (hh�eeee]r7	  (hhee]r8	  (h!]r9	  (h#h$e]r:	  (h	h�e]r;	  (hh�e]r<	  (h)heeej*	  j*	  j*	  ]r=	  (h]r>	  (h]r?	  (h]r@	  (h	h�e]rA	  (hh<e]rB	  (hhe]rC	  (h]rD	  (h	he]rE	  (hh�e]rF	  (hhe]rG	  (h]rH	  (h	he]rI	  (hh�eeee]rJ	  (hhee]rK	  (h!]rL	  (h#h$e]rM	  (h	h�e]rN	  (hh�e]rO	  (h)heee]rP	  (h]rQ	  (h]rR	  (h]rS	  (h	h�e]rT	  (hh<e]rU	  (hhe]rV	  (h]rW	  (h	he]rX	  (hh�e]rY	  (hhe]rZ	  (h]r[	  (h	he]r\	  (hh�eeee]r]	  (hhee]r^	  (h!]r_	  (h#h$e]r`	  (h	h�e]ra	  (hh�e]rb	  (h)heee]rc	  (h]rd	  (h]re	  (h]rf	  (h	h�e]rg	  (hh<e]rh	  (hhe]ri	  (h]rj	  (h	he]rk	  (hh�e]rl	  (hhe]rm	  (h]rn	  (h	he]ro	  (hh�eeee]rp	  (hhee]rq	  (h!]rr	  (h#h$e]rs	  (h	h�e]rt	  (hh�e]ru	  (h)heeejc	  ]rv	  (h]rw	  (h]rx	  (h]ry	  (h	h�e]rz	  (hh<e]r{	  (hhe]r|	  (h]r}	  (h	he]r~	  (hh�e]r	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�eeee]r�	  (hhee]r�	  (h!]r�	  (h#h$e]r�	  (h	h�e]r�	  (hh�e]r�	  (h)heeejv	  ]r�	  (h]r�	  (h]r�	  (h]r�	  (h	h�e]r�	  (hh<e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�eeee]r�	  (hhee]r�	  (h!]r�	  (h#h$e]r�	  (h	h�e]r�	  (hh�e]r�	  (h)heee]r�	  (h]r�	  (h]r�	  (h]r�	  (h	h�e]r�	  (hh<e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�eeee]r�	  (hhee]r�	  (h!]r�	  (h#h$e]r�	  (h	h�e]r�	  (hh�e]r�	  (h)heee]r�	  (h]r�	  (h]r�	  (h]r�	  (h	h
e]r�	  (hh<e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�eeee]r�	  (hhee]r�	  (h!]r�	  (h#h$e]r�	  (h	h�e]r�	  (hh�e]r�	  (h)heeej�	  ]r�	  (h]r�	  (h]r�	  (h]r�	  (h	h
e]r�	  (hh<e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�eeee]r�	  (hhee]r�	  (h!]r�	  (h#h$e]r�	  (h	h
e]r�	  (hh�e]r�	  (h)heee]r�	  (h]r�	  (h]r�	  (h]r�	  (h	h
e]r�	  (hh<e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�eeee]r�	  (hhee]r�	  (h!]r�	  (h#h$e]r�	  (h	h�e]r�	  (hh<e]r�	  (h)h�eeej�	  ]r�	  (h]r�	  (h]r�	  (h]r�	  (h	h
e]r�	  (hh<e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�e]r�	  (hhe]r�	  (h]r�	  (h	he]r�	  (hh�eeee]r�	  (hhee]r�	  (h!]r�	  (h#h$e]r�	  (h	h�e]r�	  (hh<e]r�	  (h)h�eee]r�	  (h]r�	  (h]r�	  (h]r�	  (h	h
e]r�	  (hh<e]r 
  (hhe]r
  (h]r
  (h	he]r
  (hh�e]r
  (hhe]r
  (h]r
  (h	he]r
  (hh�eeee]r
  (hhee]r	
  (h!]r

  (h#h$e]r
  (h	h
e]r
  (hh�e]r
  (h)heee]r
  (h]r
  (h]r
  (h]r
  (h	h
e]r
  (hh<e]r
  (hhe]r
  (h]r
  (h	he]r
  (hh�e]r
  (hhe]r
  (h]r
  (h	he]r
  (hh�eeee]r
  (hhee]r
  (h!]r
  (h#h$e]r
  (h	h
e]r
  (hh�e]r 
  (h)heee]r!
  (h]r"
  (h]r#
  (h]r$
  (h	h
e]r%
  (hh<e]r&
  (hhe]r'
  (h]r(
  (h	he]r)
  (hh�e]r*
  (hhe]r+
  (h]r,
  (h	he]r-
  (hh�eeee]r.
  (hhee]r/
  (h!]r0
  (h#h$e]r1
  (h	h
e]r2
  (hh�e]r3
  (h)heeej!
  ]r4
  (h]r5
  (h]r6
  (h]r7
  (h	h
e]r8
  (hh<e]r9
  (hhe]r:
  (h]r;
  (h	he]r<
  (hh�e]r=
  (hhe]r>
  (h]r?
  (h	he]r@
  (hh�eeee]rA
  (hhee]rB
  (h!]rC
  (h#h$e]rD
  (h	h
e]rE
  (hh�e]rF
  (h)heee]rG
  (h]rH
  (h]rI
  (h]rJ
  (h	h
e]rK
  (hh<e]rL
  (hhe]rM
  (h]rN
  (h	he]rO
  (hh�e]rP
  (hhe]rQ
  (h]rR
  (h	he]rS
  (hh�eeee]rT
  (hhee]rU
  (h!]rV
  (h#h$e]rW
  (h	he]rX
  (hh�e]rY
  (h)heeejG
  ]rZ
  (h]r[
  (h]r\
  (h]r]
  (h	h
e]r^
  (hh<e]r_
  (hhe]r`
  (h]ra
  (h	he]rb
  (hh�e]rc
  (hhe]rd
  (h]re
  (h	he]rf
  (hh�eeee]rg
  (hhee]rh
  (h!]ri
  (h#h$e]rj
  (h	he]rk
  (hh�e]rl
  (h)heeejZ
  jZ
  jZ
  jZ
  jZ
  ]rm
  (h]rn
  (h]ro
  (h]rp
  (h	h
e]rq
  (hh<e]rr
  (hhe]rs
  (h]rt
  (h	he]ru
  (hh�e]rv
  (hhe]rw
  (h]rx
  (h	he]ry
  (hh�eeee]rz
  (hhee]r{
  (h!]r|
  (h#h$e]r}
  (h	he]r~
  (hh�e]r
  (h)heee]r�
  (h]r�
  (h]r�
  (h]r�
  (h	h
e]r�
  (hh<e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�eeee]r�
  (hhee]r�
  (h!]r�
  (h#h$e]r�
  (h	he]r�
  (hh�e]r�
  (h)heee]r�
  (h]r�
  (h]r�
  (h]r�
  (h	h
e]r�
  (hh<e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�eeee]r�
  (hhee]r�
  (h!]r�
  (h#h$e]r�
  (h	he]r�
  (hh�e]r�
  (h)heee]r�
  (h]r�
  (h]r�
  (h]r�
  (h	h
e]r�
  (hh<e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�eeee]r�
  (hhee]r�
  (h!]r�
  (h#h$e]r�
  (h	he]r�
  (hh�e]r�
  (h)heeej�
  ]r�
  (h]r�
  (h]r�
  (h]r�
  (h	h
e]r�
  (hh<e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�eeee]r�
  (hhee]r�
  (h!]r�
  (h#h$e]r�
  (h	he]r�
  (hh�e]r�
  (h)heee]r�
  (h]r�
  (h]r�
  (h]r�
  (h	h
e]r�
  (hh<e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�eeee]r�
  (hhee]r�
  (h!]r�
  (h#h$e]r�
  (h	he]r�
  (hh�e]r�
  (h)heeej�
  ]r�
  (h]r�
  (h]r�
  (h]r�
  (h	h
e]r�
  (hh<e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�eeee]r�
  (hhee]r�
  (h!]r�
  (h#h$e]r�
  (h	he]r�
  (hh�e]r�
  (h)heeej�
  ]r�
  (h]r�
  (h]r�
  (h]r�
  (h	h
e]r�
  (hh<e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�e]r�
  (hhe]r�
  (h]r�
  (h	he]r�
  (hh�eeee]r�
  (hhee]r   (h!]r  (h#h$e]r  (h	he]r  (hh�e]r  (h)heeej�
  j�
  ]r  (h]r  (h]r  (h]r  (h	h
e]r	  (hh<e]r
  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	he]r  (hh�e]r  (h)heeej  j  j  j  j  j  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh<e]r  (hhe]r  (h]r  (h	he]r   (hh�e]r!  (hhe]r"  (h]r#  (h	he]r$  (hh�eeee]r%  (hhee]r&  (h!]r'  (h#h$e]r(  (h	he]r)  (hh�e]r*  (h)heee]r+  (h]r,  (h]r-  (h]r.  (h	h�e]r/  (hh<e]r0  (hhe]r1  (h]r2  (h	he]r3  (hh�e]r4  (hhe]r5  (h]r6  (h	he]r7  (hh�eeee]r8  (hhee]r9  (h!]r:  (h#h$e]r;  (h	j�  e]r<  (hh�e]r=  (h)heeej+  ]r>  (h]r?  (h]r@  (h]rA  (h	h�e]rB  (hh<e]rC  (hhe]rD  (h]rE  (h	he]rF  (hh�e]rG  (hhe]rH  (h]rI  (h	he]rJ  (hh�eeee]rK  (hhee]rL  (h!]rM  (h#h$e]rN  (h	j�  e]rO  (hh�e]rP  (h)heee]rQ  (h]rR  (h]rS  (h]rT  (h	h�e]rU  (hh<e]rV  (hhe]rW  (h]rX  (h	he]rY  (hh�e]rZ  (hhe]r[  (h]r\  (h	he]r]  (hh�eeee]r^  (hhee]r_  (h!]r`  (h#h$e]ra  (h	j�  e]rb  (hh�e]rc  (h)heeejQ  ]rd  (h]re  (h]rf  (h]rg  (h	h�e]rh  (hh<e]ri  (hhe]rj  (h]rk  (h	he]rl  (hh�e]rm  (hhe]rn  (h]ro  (h	he]rp  (hh�eeee]rq  (hhee]rr  (h!]rs  (h#h$e]rt  (h	j�  e]ru  (hh<e]rv  (h)heee]rw  (h]rx  (h]ry  (h]rz  (h	h�e]r{  (hh<e]r|  (hhe]r}  (h]r~  (h	he]r  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)heeejw  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r   (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�eeee]r	  (hhee]r
  (h!]r  (h#h$e]r  (h	he]r  (hh<e]r  (h)heee]r  (h]r  (h]r  (h]r  (h	h
e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	he]r   (hh<e]r!  (h)heeej  j  j  j  j  j  ]r"  (h]r#  (h]r$  (h]r%  (h	h
e]r&  (hh�e]r'  (hhe]r(  (h]r)  (h	he]r*  (hh�e]r+  (hhe]r,  (h]r-  (h	he]r.  (hh�eeee]r/  (hhee]r0  (h!]r1  (h#h$e]r2  (h	he]r3  (hh<e]r4  (h)heee]r5  (h]r6  (h]r7  (h]r8  (h	h
e]r9  (hh�e]r:  (hhe]r;  (h]r<  (h	he]r=  (hh�e]r>  (hhe]r?  (h]r@  (h	he]rA  (hh�eeee]rB  (hhee]rC  (h!]rD  (h#h$e]rE  (h	he]rF  (hh<e]rG  (h)heeej5  j5  j5  j5  ]rH  (h]rI  (h]rJ  (h]rK  (h	h
e]rL  (hh�e]rM  (hhe]rN  (h]rO  (h	h�e]rP  (hh�e]rQ  (hhe]rR  (h]rS  (h	he]rT  (hh�eeee]rU  (hhee]rV  (h!]rW  (h#h$e]rX  (h	he]rY  (hh<e]rZ  (h)heee]r[  (h]r\  (h]r]  (h]r^  (h	h
e]r_  (hh�e]r`  (hhe]ra  (h]rb  (h	h�e]rc  (hh�e]rd  (hhe]re  (h]rf  (h	he]rg  (hh�eeee]rh  (hhee]ri  (h!]rj  (h#h$e]rk  (h	j�  e]rl  (hh�e]rm  (h)h�eee]rn  (h]ro  (h]rp  (h]rq  (h	h
e]rr  (hh�e]rs  (hhe]rt  (h]ru  (h	h�e]rv  (hh�e]rw  (hhe]rx  (h]ry  (h	he]rz  (hh�eeee]r{  (hhee]r|  (h!]r}  (h#h$e]r~  (h	j�  e]r  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�eeee]r   (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)h�eeej�  j�  j�  j�  j�  j�  j�  j�  ]r  (h]r  (h]r  (h]r	  (h	h
e]r
  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)h�eeej  j  ]r  (h]r  (h]r  (h]r  (h	h
e]r  (hh�e]r  (hhe]r  (h]r   (h	he]r!  (hh�e]r"  (hhe]r#  (h]r$  (h	he]r%  (hh�eeee]r&  (hhee]r'  (h!]r(  (h#h$e]r)  (h	j�  e]r*  (hh�e]r+  (h)h�eeej  j  j  ]r,  (h]r-  (h]r.  (h]r/  (h	h
e]r0  (hh�e]r1  (hhe]r2  (h]r3  (h	he]r4  (hh�e]r5  (hhe]r6  (h]r7  (h	he]r8  (hh�eeee]r9  (hhee]r:  (h!]r;  (h#h$e]r<  (h	j�  e]r=  (hh�e]r>  (h)h�eee]r?  (h]r@  (h]rA  (h]rB  (h	h
e]rC  (hh�e]rD  (hhe]rE  (h]rF  (h	he]rG  (hh�e]rH  (hhe]rI  (h]rJ  (h	he]rK  (hh�eeee]rL  (hhee]rM  (h!]rN  (h#h$e]rO  (h	j�  e]rP  (hh�e]rQ  (h)h�eee]rR  (h]rS  (h]rT  (h]rU  (h	h
e]rV  (hh�e]rW  (hhe]rX  (h]rY  (h	he]rZ  (hh�e]r[  (hhe]r\  (h]r]  (h	he]r^  (hh�eeee]r_  (hhee]r`  (h!]ra  (h#h$e]rb  (h	j�  e]rc  (hh�e]rd  (h)h�eee]re  (h]rf  (h]rg  (h]rh  (h	h
e]ri  (hh�e]rj  (hhe]rk  (h]rl  (h	he]rm  (hh�e]rn  (hhe]ro  (h]rp  (h	he]rq  (hh�eeee]rr  (hhee]rs  (h!]rt  (h#h$e]ru  (h	h
e]rv  (hh�e]rw  (h)h�eee]rx  (h]ry  (h]rz  (h]r{  (h	h
e]r|  (hh�e]r}  (hhe]r~  (h]r  (h	he]r�  (hh�e]r�  (hhe]r�  (X	   Next-Mover�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r   (h]r  (h	h
e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (j�  ]r	  (h	he]r
  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	h
e]r  (hh�e]r  (h)heeej�  ]r  (h]r  (h]r  (h]r  (h	h
e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (j�  ]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r   (h#h$e]r!  (h	h
e]r"  (hh�e]r#  (h)heee]r$  (h]r%  (h]r&  (h]r'  (h	h
e]r(  (hh�e]r)  (hhe]r*  (h]r+  (h	he]r,  (hh�e]r-  (hhe]r.  (j�  ]r/  (h	he]r0  (hh�eeee]r1  (hhee]r2  (h!]r3  (h#h$e]r4  (h	j�  e]r5  (hh�e]r6  (h)heee]r7  (h]r8  (h]r9  (h]r:  (h	h
e]r;  (hh�e]r<  (hhe]r=  (h]r>  (h	he]r?  (hh�e]r@  (hhe]rA  (j�  ]rB  (h	he]rC  (hh�eeee]rD  (hhee]rE  (h!]rF  (h#h$e]rG  (h	j�  e]rH  (hh�e]rI  (h)heee]rJ  (h]rK  (h]rL  (h]rM  (h	h
e]rN  (hh�e]rO  (hhe]rP  (h]rQ  (h	he]rR  (hh�e]rS  (hhe]rT  (j�  ]rU  (h	he]rV  (hh�eeee]rW  (hhee]rX  (h!]rY  (h#h$e]rZ  (h	he]r[  (hh<e]r\  (h)h�eee]r]  (h]r^  (h]r_  (h]r`  (h	h
e]ra  (hh�e]rb  (hhe]rc  (h]rd  (h	h�e]re  (hh�e]rf  (hhe]rg  (j�  ]rh  (h	he]ri  (hh�eeee]rj  (hhee]rk  (h!]rl  (h#h$e]rm  (h	he]rn  (hh<e]ro  (h)h�eeej]  ]rp  (h]rq  (h]rr  (h]rs  (h	h
e]rt  (hh�e]ru  (hhe]rv  (h]rw  (h	h�e]rx  (hh�e]ry  (hhe]rz  (j�  ]r{  (h	he]r|  (hh�eeee]r}  (hhee]r~  (h!]r  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)h�eeejp  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (X	   Next-Mover�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)h�eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)h�eeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)h�eeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)h�eee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)h�eeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r   (j�  ]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	h�e]r  (hh�e]r  (h)h�eeej�  ]r	  (h]r
  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	h�e]r  (hh�e]r  (h)heee]r  (h]r  (h]r  (h]r  (h	h�e]r   (hh�e]r!  (hhe]r"  (h]r#  (h	h�e]r$  (hh�e]r%  (hhe]r&  (j�  ]r'  (h	he]r(  (hh�eeee]r)  (hhee]r*  (h!]r+  (h#h$e]r,  (h	h�e]r-  (hh�e]r.  (h)heee]r/  (h]r0  (h]r1  (h]r2  (h	h�e]r3  (hh�e]r4  (hhe]r5  (h]r6  (h	h�e]r7  (hh�e]r8  (hhe]r9  (j�  ]r:  (h	he]r;  (hh�eeee]r<  (hhee]r=  (h!]r>  (h#h$e]r?  (h	h�e]r@  (hh�e]rA  (h)heeej/  j/  j/  j/  ]rB  (h]rC  (h]rD  (h]rE  (h	h�e]rF  (hh�e]rG  (hhe]rH  (h]rI  (h	h�e]rJ  (hh�e]rK  (hhe]rL  (j�  ]rM  (h	he]rN  (hh�eeee]rO  (hhee]rP  (h!]rQ  (h#h$e]rR  (h	h�e]rS  (hh�e]rT  (h)heeejB  jB  jB  ]rU  (h]rV  (h]rW  (h]rX  (h	h�e]rY  (hh�e]rZ  (hhe]r[  (h]r\  (h	h�e]r]  (hh�e]r^  (hhe]r_  (j�  ]r`  (h	he]ra  (hh�eeee]rb  (hhee]rc  (h!]rd  (h#h$e]re  (h	h�e]rf  (hh�e]rg  (h)heeejU  jU  jU  ]rh  (h]ri  (h]rj  (h]rk  (h	h�e]rl  (hh�e]rm  (hhe]rn  (h]ro  (h	h�e]rp  (hh�e]rq  (hhe]rr  (j�  ]rs  (h	he]rt  (hh�eeee]ru  (hhee]rv  (h!]rw  (h#h$e]rx  (h	h�e]ry  (hh�e]rz  (h)heee]r{  (h]r|  (h]r}  (h]r~  (h	h�e]r  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)heeej{  j{  j{  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)h�eee]r   (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r	  (hhe]r
  (j�  ]r  (h	he]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh<e]r  (h)h�eee]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	he]r  (hh�eeee]r   (hhee]r!  (h!]r"  (h#h$e]r#  (h	j�  e]r$  (hh<e]r%  (h)h�eee]r&  (h]r'  (h]r(  (h]r)  (h	h�e]r*  (hh�e]r+  (hhe]r,  (h]r-  (h	h�e]r.  (hh�e]r/  (hhe]r0  (j�  ]r1  (h	he]r2  (hh�eeee]r3  (hhee]r4  (h!]r5  (h#h$e]r6  (h	j�  e]r7  (hh<e]r8  (h)h�eeej&  ]r9  (h]r:  (h]r;  (h]r<  (h	h�e]r=  (hh�e]r>  (hhe]r?  (h]r@  (h	h�e]rA  (hh�e]rB  (hhe]rC  (j�  ]rD  (h	he]rE  (hh�eeee]rF  (hhee]rG  (h!]rH  (h#h$e]rI  (h	j�  e]rJ  (hh�e]rK  (h)h�eeej9  ]rL  (h]rM  (h]rN  (h]rO  (h	h�e]rP  (hh�e]rQ  (hhe]rR  (h]rS  (h	h�e]rT  (hh�e]rU  (hhe]rV  (j�  ]rW  (h	h�e]rX  (hh�eeee]rY  (hhee]rZ  (h!]r[  (h#h$e]r\  (h	j�  e]r]  (hh�e]r^  (h)h�eee]r_  (h]r`  (h]ra  (h]rb  (h	h�e]rc  (hh�e]rd  (hhe]re  (h]rf  (h	h�e]rg  (hh�e]rh  (hhe]ri  (j�  ]rj  (h	h�e]rk  (hh�eeee]rl  (hhee]rm  (h!]rn  (h#h$e]ro  (h	j�  e]rp  (hh�e]rq  (h)h�eeej_  ]rr  (h]rs  (h]rt  (h]ru  (h	h�e]rv  (hh�e]rw  (hhe]rx  (h]ry  (h	h�e]rz  (hh�e]r{  (hhe]r|  (j�  ]r}  (h	h�e]r~  (hh�eeee]r  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)h�eeejr  jr  jr  jr  jr  jr  jr  jr  jr  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r   (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r	  (h)heeej�  ]r
  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej
  j
  j
  j
  ]r  (h]r  (h]r  (h]r   (h	h�e]r!  (hh�e]r"  (hhe]r#  (h]r$  (h	h�e]r%  (hh�e]r&  (hhe]r'  (j�  ]r(  (h	h�e]r)  (hh�eeee]r*  (hhee]r+  (h!]r,  (h#h$e]r-  (h	j�  e]r.  (hh�e]r/  (h)heeej  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  j  ]r0  (h]r1  (h]r2  (h]r3  (h	h�e]r4  (hh�e]r5  (hhe]r6  (h]r7  (h	h�e]r8  (hh�e]r9  (hhe]r:  (j�  ]r;  (h	h�e]r<  (hh�eeee]r=  (hhee]r>  (h!]r?  (h#h$e]r@  (h	j�  e]rA  (hh�e]rB  (h)heeej0  j0  j0  j0  j0  j0  j0  ]rC  (h]rD  (h]rE  (h]rF  (h	h�e]rG  (hh�e]rH  (hhe]rI  (h]rJ  (h	he]rK  (hh�e]rL  (hhe]rM  (j�  ]rN  (h	h�e]rO  (hh�eeee]rP  (hhee]rQ  (h!]rR  (h#h$e]rS  (h	j�  e]rT  (hh�e]rU  (h)heeejC  ]rV  (h]rW  (h]rX  (h]rY  (h	h�e]rZ  (hh�e]r[  (hhe]r\  (h]r]  (h	he]r^  (hh�e]r_  (hhe]r`  (j�  ]ra  (h	h�e]rb  (hh�eeee]rc  (hhee]rd  (h!]re  (h#h$e]rf  (h	j�  e]rg  (hh�e]rh  (h)heee]ri  (h]rj  (h]rk  (h]rl  (h	h�e]rm  (hh�e]rn  (hhe]ro  (h]rp  (h	he]rq  (hh�e]rr  (hhe]rs  (j�  ]rt  (h	h�e]ru  (hh�eeee]rv  (hhee]rw  (h!]rx  (h#h$e]ry  (h	j�  e]rz  (hh�e]r{  (h)heeeji  ji  ji  ]r|  (h]r}  (h]r~  (h]r  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej|  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r   (h)heeej�  j�  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r	  (hh�e]r
  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej  j  j  j  j  j  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r   (hh�eeee]r!  (hhee]r"  (h!]r#  (h#h$e]r$  (h	j�  e]r%  (hh�e]r&  (h)heeej  ]r'  (h]r(  (h]r)  (h]r*  (h	h�e]r+  (hh�e]r,  (hhe]r-  (h]r.  (h	he]r/  (hh�e]r0  (hhe]r1  (j�  ]r2  (h	h�e]r3  (hh�eeee]r4  (hhee]r5  (h!]r6  (h#h$e]r7  (h	j�  e]r8  (hh�e]r9  (h)heeej'  j'  j'  j'  j'  j'  j'  ]r:  (h]r;  (h]r<  (h]r=  (h	h�e]r>  (hh�e]r?  (hhe]r@  (h]rA  (h	he]rB  (hh�e]rC  (hhe]rD  (j�  ]rE  (h	h�e]rF  (hh�eeee]rG  (hhee]rH  (h!]rI  (h#h$e]rJ  (h	j�  e]rK  (hh�e]rL  (h)heeej:  j:  j:  j:  j:  j:  j:  ]rM  (h]rN  (h]rO  (h]rP  (h	h�e]rQ  (hh�e]rR  (hhe]rS  (h]rT  (h	he]rU  (hh�e]rV  (hhe]rW  (j�  ]rX  (h	h�e]rY  (hh�eeee]rZ  (hhee]r[  (h!]r\  (h#h$e]r]  (h	j�  e]r^  (hh�e]r_  (h)heeejM  ]r`  (h]ra  (h]rb  (h]rc  (h	h�e]rd  (hh�e]re  (hhe]rf  (h]rg  (h	h�e]rh  (hh�e]ri  (hhe]rj  (j�  ]rk  (h	h�e]rl  (hh�eeee]rm  (hhee]rn  (h!]ro  (h#h$e]rp  (h	j�  e]rq  (hh�e]rr  (h)heee]rs  (h]rt  (h]ru  (h]rv  (h	h�e]rw  (hh�e]rx  (hhe]ry  (h]rz  (h	h�e]r{  (hh�e]r|  (hhe]r}  (j�  ]r~  (h	h�e]r  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeejs  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r   (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r	  (hh�e]r
  (h)heee]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heee]r  (h]r  (h]r   (h]r!  (h	h�e]r"  (hh�e]r#  (hhe]r$  (h]r%  (h	he]r&  (hh�e]r'  (hhe]r(  (j�  ]r)  (h	h�e]r*  (hh�eeee]r+  (hhee]r,  (h!]r-  (h#h$e]r.  (h	j�  e]r/  (hh�e]r0  (h)heeej  ]r1  (h]r2  (h]r3  (h]r4  (h	h�e]r5  (hh�e]r6  (hhe]r7  (h]r8  (h	he]r9  (hh�e]r:  (hhe]r;  (j�  ]r<  (h	h�e]r=  (hh�eeee]r>  (hhee]r?  (h!]r@  (h#h$e]rA  (h	j�  e]rB  (hh�e]rC  (h)heeej1  j1  ]rD  (h]rE  (h]rF  (h]rG  (h	h�e]rH  (hh�e]rI  (hhe]rJ  (h]rK  (h	he]rL  (hh�e]rM  (hhe]rN  (j�  ]rO  (h	h�e]rP  (hh�eeee]rQ  (hhee]rR  (h!]rS  (h#h$e]rT  (h	j�  e]rU  (hh�e]rV  (h)heeejD  jD  jD  jD  jD  jD  jD  jD  jD  jD  ]rW  (h]rX  (h]rY  (h]rZ  (h	h�e]r[  (hh�e]r\  (hhe]r]  (h]r^  (h	he]r_  (hh�e]r`  (hhe]ra  (j�  ]rb  (h	h�e]rc  (hh�eeee]rd  (hhee]re  (h!]rf  (h#h$e]rg  (h	j�  e]rh  (hh�e]ri  (h)heeejW  jW  jW  jW  jW  jW  ]rj  (h]rk  (h]rl  (h]rm  (h	h�e]rn  (hh�e]ro  (hhe]rp  (h]rq  (h	he]rr  (hh�e]rs  (hhe]rt  (j�  ]ru  (h	h�e]rv  (hh�eeee]rw  (hhee]rx  (h!]ry  (h#h$e]rz  (h	j�  e]r{  (hh�e]r|  (h)heee]r}  (h]r~  (h]r  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (X	   Next-Mover�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r   (h	j�  e]r  (hh�e]r  (h)heeej�  j�  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r	  (h]r
  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej  j  j  j  j  j  j  j  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r   (j�  ]r!  (h	h�e]r"  (hh�eeee]r#  (hhee]r$  (h!]r%  (h#h$e]r&  (h	j�  e]r'  (hh�e]r(  (h)heeej  j  ]r)  (h]r*  (h]r+  (h]r,  (h	h�e]r-  (hh�e]r.  (hhe]r/  (h]r0  (h	h�e]r1  (hh�e]r2  (hhe]r3  (j�  ]r4  (h	h�e]r5  (hh�eeee]r6  (hhee]r7  (h!]r8  (h#h$e]r9  (h	j�  e]r:  (hh�e]r;  (h)heeej)  j)  j)  j)  ]r<  (h]r=  (h]r>  (h]r?  (h	h�e]r@  (hh�e]rA  (hhe]rB  (h]rC  (h	h�e]rD  (hh�e]rE  (hhe]rF  (j�  ]rG  (h	h�e]rH  (hh�eeee]rI  (hhee]rJ  (h!]rK  (h#h$e]rL  (h	j�  e]rM  (hh�e]rN  (h)heeej<  j<  ]rO  (h]rP  (h]rQ  (h]rR  (h	h�e]rS  (hh�e]rT  (hhe]rU  (h]rV  (h	h�e]rW  (hh�e]rX  (hhe]rY  (j�  ]rZ  (h	h�e]r[  (hh�eeee]r\  (hhee]r]  (h!]r^  (h#h$e]r_  (h	j�  e]r`  (hh�e]ra  (h)heeejO  ]rb  (h]rc  (h]rd  (h]re  (h	h�e]rf  (hh�e]rg  (hhe]rh  (h]ri  (h	h�e]rj  (hh�e]rk  (hhe]rl  (j�  ]rm  (h	h�e]rn  (hh�eeee]ro  (hhee]rp  (h!]rq  (h#h$e]rr  (h	j�  e]rs  (hh�e]rt  (h)heeejb  ]ru  (h]rv  (h]rw  (h]rx  (h	h�e]ry  (hh�e]rz  (hhe]r{  (h]r|  (h	h�e]r}  (hh�e]r~  (hhe]r  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeeju  ju  ju  ju  ju  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r   (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r	  (h#h$e]r
  (h	j�  e]r  (hh�e]r  (h)heee]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heee]r   (h]r!  (h]r"  (h]r#  (h	h�e]r$  (hh�e]r%  (hhe]r&  (h]r'  (h	he]r(  (hh�e]r)  (hhe]r*  (j�  ]r+  (h	h�e]r,  (hh�eeee]r-  (hhee]r.  (h!]r/  (h#h$e]r0  (h	j�  e]r1  (hh�e]r2  (h)heeej   j   j   j   ]r3  (h]r4  (h]r5  (h]r6  (h	h�e]r7  (hh�e]r8  (hhe]r9  (h]r:  (h	he]r;  (hh�e]r<  (hhe]r=  (j�  ]r>  (h	h�e]r?  (hh�eeee]r@  (hhee]rA  (h!]rB  (h#h$e]rC  (h	j�  e]rD  (hh�e]rE  (h)heeej3  j3  j3  j3  j3  j3  j3  ]rF  (h]rG  (h]rH  (h]rI  (h	h�e]rJ  (hh�e]rK  (hhe]rL  (h]rM  (h	he]rN  (hh�e]rO  (hhe]rP  (j�  ]rQ  (h	h�e]rR  (hh�eeee]rS  (hhee]rT  (h!]rU  (h#h$e]rV  (h	j�  e]rW  (hh�e]rX  (h)heeejF  ]rY  (h]rZ  (h]r[  (h]r\  (h	h�e]r]  (hh�e]r^  (hhe]r_  (h]r`  (h	he]ra  (hh�e]rb  (hhe]rc  (j�  ]rd  (h	h�e]re  (hh�eeee]rf  (hhee]rg  (h!]rh  (h#h$e]ri  (h	j�  e]rj  (hh�e]rk  (h)heeejY  jY  jY  jY  jY  jY  ]rl  (h]rm  (h]rn  (h]ro  (h	h�e]rp  (hh�e]rq  (hhe]rr  (h]rs  (h	he]rt  (hh�e]ru  (hhe]rv  (j�  ]rw  (h	h�e]rx  (hh�eeee]ry  (hhee]rz  (h!]r{  (h#h$e]r|  (h	j�  e]r}  (hh�e]r~  (h)heeejl  jl  ]r  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej  j  j  j  j  j  j  j  j  j  j  j  j  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r   (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej�  j�  j�  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r	  (hhe]r
  (h]r  (h	he]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r   (hhe]r!  (j�  ]r"  (h	h�e]r#  (hh�eeee]r$  (hhee]r%  (h!]r&  (h#h$e]r'  (h	j�  e]r(  (hh�e]r)  (h)heeej  j  j  j  ]r*  (h]r+  (h]r,  (h]r-  (h	h�e]r.  (hh�e]r/  (hhe]r0  (h]r1  (h	he]r2  (hh�e]r3  (hhe]r4  (j�  ]r5  (h	h�e]r6  (hh�eeee]r7  (hhee]r8  (h!]r9  (h#h$e]r:  (h	j�  e]r;  (hh�e]r<  (h)heee]r=  (h]r>  (h]r?  (h]r@  (h	h�e]rA  (hh�e]rB  (hhe]rC  (h]rD  (h	h�e]rE  (hh�e]rF  (hhe]rG  (j�  ]rH  (h	h�e]rI  (hh�eeee]rJ  (hhee]rK  (h!]rL  (h#h$e]rM  (h	j�  e]rN  (hh�e]rO  (h)heee]rP  (h]rQ  (h]rR  (h]rS  (h	h�e]rT  (hh�e]rU  (hhe]rV  (h]rW  (h	h�e]rX  (hh�e]rY  (hhe]rZ  (j�  ]r[  (h	h�e]r\  (hh�eeee]r]  (hhee]r^  (h!]r_  (h#h$e]r`  (h	j�  e]ra  (hh�e]rb  (h)heeejP  jP  jP  jP  jP  jP  ]rc  (h]rd  (h]re  (h]rf  (h	h�e]rg  (hh�e]rh  (hhe]ri  (h]rj  (h	h�e]rk  (hh�e]rl  (hhe]rm  (j�  ]rn  (h	h�e]ro  (hh�eeee]rp  (hhee]rq  (h!]rr  (h#h$e]rs  (h	j�  e]rt  (hh�e]ru  (h)heeejc  jc  jc  ]rv  (h]rw  (h]rx  (h]ry  (h	h�e]rz  (hh�e]r{  (hhe]r|  (h]r}  (h	h�e]r~  (hh�e]r  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeejv  jv  jv  jv  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r   (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r	  (h!]r
  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heee]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r   (h)heeej  j  ]r!  (h]r"  (h]r#  (h]r$  (h	h�e]r%  (hh�e]r&  (hhe]r'  (h]r(  (h	h�e]r)  (hh�e]r*  (hhe]r+  (j�  ]r,  (h	h�e]r-  (hh�eeee]r.  (hhee]r/  (h!]r0  (h#h$e]r1  (h	j�  e]r2  (hh�e]r3  (h)heeej!  j!  ]r4  (h]r5  (h]r6  (h]r7  (h	h�e]r8  (hh�e]r9  (hhe]r:  (h]r;  (h	h�e]r<  (hh�e]r=  (hhe]r>  (j�  ]r?  (h	h�e]r@  (hh�eeee]rA  (hhee]rB  (h!]rC  (h#h$e]rD  (h	j�  e]rE  (hh�e]rF  (h)heee]rG  (h]rH  (h]rI  (h]rJ  (h	h�e]rK  (hh�e]rL  (hhe]rM  (h]rN  (h	h�e]rO  (hh�e]rP  (hhe]rQ  (j�  ]rR  (h	h�e]rS  (hh�eeee]rT  (hhee]rU  (h!]rV  (h#h$e]rW  (h	j�  e]rX  (hh�e]rY  (h)heeejG  jG  jG  jG  jG  jG  jG  jG  jG  jG  jG  ]rZ  (h]r[  (h]r\  (h]r]  (h	h�e]r^  (hh�e]r_  (hhe]r`  (h]ra  (h	h�e]rb  (hh�e]rc  (hhe]rd  (j�  ]re  (h	h�e]rf  (hh�eeee]rg  (hhee]rh  (h!]ri  (h#h$e]rj  (h	j�  e]rk  (hh�e]rl  (h)heee]rm  (h]rn  (h]ro  (h]rp  (h	h�e]rq  (hh�e]rr  (hhe]rs  (h]rt  (h	h�e]ru  (hh�e]rv  (hhe]rw  (j�  ]rx  (h	h�e]ry  (hh�eeee]rz  (hhee]r{  (h!]r|  (h#h$e]r}  (h	j�  e]r~  (hh�e]r  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r   (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej�  ]r  (h]r  (h]r  (h]r  (h	h�e]r	  (hh�e]r
  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r   (hh�e]r!  (hhe]r"  (j�  ]r#  (h	h�e]r$  (hh�eeee]r%  (hhee]r&  (h!]r'  (h#h$e]r(  (h	j�  e]r)  (hh�e]r*  (h)heeej  j  j  j  ]r+  (h]r,  (h]r-  (h]r.  (h	h�e]r/  (hh�e]r0  (hhe]r1  (h]r2  (h	h�e]r3  (hh�e]r4  (hhe]r5  (j�  ]r6  (h	h�e]r7  (hh�eeee]r8  (hhee]r9  (h!]r:  (h#h$e]r;  (h	j�  e]r<  (hh�e]r=  (h)heeej+  j+  j+  j+  j+  ]r>  (h]r?  (h]r@  (h]rA  (h	h�e]rB  (hh�e]rC  (hhe]rD  (h]rE  (h	h�e]rF  (hh�e]rG  (hhe]rH  (j�  ]rI  (h	h�e]rJ  (hh�eeee]rK  (hhee]rL  (h!]rM  (h#h$e]rN  (h	j�  e]rO  (hh�e]rP  (h)heee]rQ  (h]rR  (h]rS  (h]rT  (h	h�e]rU  (hh�e]rV  (hhe]rW  (h]rX  (h	h�e]rY  (hh�e]rZ  (hhe]r[  (j�  ]r\  (h	h�e]r]  (hh�eeee]r^  (hhee]r_  (h!]r`  (h#h$e]ra  (h	j�  e]rb  (hh�e]rc  (h)heeejQ  jQ  jQ  jQ  ]rd  (h]re  (h]rf  (h]rg  (h	h�e]rh  (hh�e]ri  (hhe]rj  (h]rk  (h	h�e]rl  (hh�e]rm  (hhe]rn  (j�  ]ro  (h	h�e]rp  (hh�eeee]rq  (hhee]rr  (h!]rs  (h#h$e]rt  (h	j�  e]ru  (hh�e]rv  (h)heeejd  jd  jd  jd  ]rw  (h]rx  (h]ry  (h]rz  (h	h�e]r{  (hh�e]r|  (hhe]r}  (h]r~  (h	h�e]r  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r   (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r	  (hhee]r
  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r   (hh�e]r!  (h)heeej  j  j  j  ]r"  (h]r#  (h]r$  (h]r%  (h	h�e]r&  (hh�e]r'  (hhe]r(  (h]r)  (h	he]r*  (hh�e]r+  (hhe]r,  (j�  ]r-  (h	h�e]r.  (hh�eeee]r/  (hhee]r0  (h!]r1  (h#h$e]r2  (h	j�  e]r3  (hh�e]r4  (h)heee]r5  (h]r6  (h]r7  (h]r8  (h	h�e]r9  (hh�e]r:  (hhe]r;  (h]r<  (h	he]r=  (hh�e]r>  (hhe]r?  (j�  ]r@  (h	h�e]rA  (hh�eeee]rB  (hhee]rC  (h!]rD  (h#h$e]rE  (h	j�  e]rF  (hh�e]rG  (h)heee]rH  (h]rI  (h]rJ  (h]rK  (h	h�e]rL  (hh�e]rM  (hhe]rN  (h]rO  (h	he]rP  (hh�e]rQ  (hhe]rR  (j�  ]rS  (h	h�e]rT  (hh�eeee]rU  (hhee]rV  (h!]rW  (h#h$e]rX  (h	j�  e]rY  (hh�e]rZ  (h)heee]r[  (h]r\  (h]r]  (h]r^  (h	h�e]r_  (hh�e]r`  (hhe]ra  (h]rb  (h	he]rc  (hh�e]rd  (hhe]re  (j�  ]rf  (h	h�e]rg  (hh�eeee]rh  (hhee]ri  (h!]rj  (h#h$e]rk  (h	j�  e]rl  (hh�e]rm  (h)heeej[  ]rn  (h]ro  (h]rp  (h]rq  (h	h�e]rr  (hh�e]rs  (hhe]rt  (h]ru  (h	he]rv  (hh�e]rw  (hhe]rx  (j�  ]ry  (h	h�e]rz  (hh�eeee]r{  (hhee]r|  (h!]r}  (h#h$e]r~  (h	j�  e]r  (hh�e]r�  (h)heeejn  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r   (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej�  j�  j�  j�  j�  j�  j�  ]r  (h]r  (h]r  (h]r	  (h	h�e]r
  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heee]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r   (h	he]r!  (hh�e]r"  (hhe]r#  (j�  ]r$  (h	h�e]r%  (hh�eeee]r&  (hhee]r'  (h!]r(  (h#h$e]r)  (h	j�  e]r*  (hh�e]r+  (h)heeej  ]r,  (h]r-  (h]r.  (h]r/  (h	h�e]r0  (hh�e]r1  (hhe]r2  (h]r3  (h	he]r4  (hh�e]r5  (hhe]r6  (j�  ]r7  (h	h�e]r8  (hh�eeee]r9  (hhee]r:  (h!]r;  (h#h$e]r<  (h	j�  e]r=  (hh�e]r>  (h)heeej,  j,  j,  j,  j,  j,  j,  j,  ]r?  (h]r@  (h]rA  (h]rB  (h	h�e]rC  (hh�e]rD  (hhe]rE  (h]rF  (h	he]rG  (hh�e]rH  (hhe]rI  (j�  ]rJ  (h	h�e]rK  (hh�eeee]rL  (hhee]rM  (h!]rN  (h#h$e]rO  (h	j�  e]rP  (hh�e]rQ  (h)heee]rR  (h]rS  (h]rT  (h]rU  (h	h�e]rV  (hh�e]rW  (hhe]rX  (h]rY  (h	he]rZ  (hh�e]r[  (hhe]r\  (j�  ]r]  (h	h�e]r^  (hh�eeee]r_  (hhee]r`  (h!]ra  (h#h$e]rb  (h	j�  e]rc  (hh�e]rd  (h)heeejR  jR  ]re  (h]rf  (h]rg  (h]rh  (h	h�e]ri  (hh�e]rj  (hhe]rk  (h]rl  (h	he]rm  (hh�e]rn  (hhe]ro  (j�  ]rp  (h	h�e]rq  (hh�eeee]rr  (hhee]rs  (h!]rt  (h#h$e]ru  (h	j�  e]rv  (hh�e]rw  (h)heeeje  ]rx  (h]ry  (h]rz  (h]r{  (h	h�e]r|  (hh�e]r}  (hhe]r~  (h]r  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeejx  e(jx  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r   (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r	  (hh�eeee]r
  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej�  j�  j�  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r   (h	j�  e]r!  (hh�e]r"  (h)heeej  ]r#  (h]r$  (h]r%  (h]r&  (h	h�e]r'  (hh�e]r(  (hhe]r)  (h]r*  (h	h�e]r+  (hh�e]r,  (hhe]r-  (j�  ]r.  (h	h�e]r/  (hh�eeee]r0  (hhee]r1  (h!]r2  (h#h$e]r3  (h	j�  e]r4  (hh�e]r5  (h)heee]r6  (h]r7  (h]r8  (h]r9  (h	h�e]r:  (hh�e]r;  (hhe]r<  (h]r=  (h	h�e]r>  (hh�e]r?  (hhe]r@  (j�  ]rA  (h	h�e]rB  (hh�eeee]rC  (hhee]rD  (h!]rE  (h#h$e]rF  (h	j�  e]rG  (hh�e]rH  (h)heee]rI  (h]rJ  (h]rK  (h]rL  (h	h�e]rM  (hh�e]rN  (hhe]rO  (h]rP  (h	h�e]rQ  (hh�e]rR  (hhe]rS  (j�  ]rT  (h	h�e]rU  (hh�eeee]rV  (hhee]rW  (h!]rX  (h#h$e]rY  (h	j�  e]rZ  (hh�e]r[  (h)heeejI  jI  ]r\  (h]r]  (h]r^  (h]r_  (h	h�e]r`  (hh�e]ra  (hhe]rb  (h]rc  (h	h�e]rd  (hh�e]re  (hhe]rf  (j�  ]rg  (h	h�e]rh  (hh�eeee]ri  (hhee]rj  (h!]rk  (h#h$e]rl  (h	j�  e]rm  (hh�e]rn  (h)heeej\  j\  j\  j\  ]ro  (h]rp  (h]rq  (h]rr  (h	h�e]rs  (hh�e]rt  (hhe]ru  (h]rv  (h	h�e]rw  (hh�e]rx  (hhe]ry  (j�  ]rz  (h	h�e]r{  (hh�eeee]r|  (hhee]r}  (h!]r~  (h#h$e]r  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r   (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heee]r  (h]r  (h]r	  (h]r
  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej  j  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r   (h]r!  (h	h�e]r"  (hh�e]r#  (hhe]r$  (j�  ]r%  (h	h�e]r&  (hh�eeee]r'  (hhee]r(  (h!]r)  (h#h$e]r*  (h	j�  e]r+  (hh�e]r,  (h)heeej  j  j  ]r-  (h]r.  (h]r/  (h]r0  (h	h�e]r1  (hh�e]r2  (hhe]r3  (h]r4  (h	h�e]r5  (hh�e]r6  (hhe]r7  (j�  ]r8  (h	h�e]r9  (hh�eeee]r:  (hhee]r;  (h!]r<  (h#h$e]r=  (h	j�  e]r>  (hh�e]r?  (h)heeej-  j-  j-  j-  j-  j-  j-  j-  j-  j-  ]r@  (h]rA  (h]rB  (h]rC  (h	h�e]rD  (hh�e]rE  (hhe]rF  (h]rG  (h	h�e]rH  (hh�e]rI  (hhe]rJ  (j�  ]rK  (h	h�e]rL  (hh�eeee]rM  (hhee]rN  (h!]rO  (h#h$e]rP  (h	j�  e]rQ  (hh�e]rR  (h)heee]rS  (h]rT  (h]rU  (h]rV  (h	h�e]rW  (hh�e]rX  (hhe]rY  (h]rZ  (h	h�e]r[  (hh�e]r\  (hhe]r]  (j�  ]r^  (h	h�e]r_  (hh�eeee]r`  (hhee]ra  (h!]rb  (h#h$e]rc  (h	j�  e]rd  (hh�e]re  (h)heeejS  ]rf  (h]rg  (h]rh  (h]ri  (h	h�e]rj  (hh�e]rk  (hhe]rl  (h]rm  (h	h�e]rn  (hh�e]ro  (hhe]rp  (j�  ]rq  (h	h�e]rr  (hh�eeee]rs  (hhee]rt  (h!]ru  (h#h$e]rv  (h	j�  e]rw  (hh�e]rx  (h)heeejf  ]ry  (h]rz  (h]r{  (h]r|  (h	h�e]r}  (hh�e]r~  (hhe]r  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeejy  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r   (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r	  (h	h�e]r
  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heee]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r   (h#h$e]r!  (h	j�  e]r"  (hh�e]r#  (h)heeej  j  j  j  j  j  j  ]r$  (h]r%  (h]r&  (h]r'  (h	h�e]r(  (hh�e]r)  (hhe]r*  (h]r+  (h	h�e]r,  (hh�e]r-  (hhe]r.  (j�  ]r/  (h	h�e]r0  (hh�eeee]r1  (hhee]r2  (h!]r3  (h#h$e]r4  (h	j�  e]r5  (hh�e]r6  (h)heeej$  ]r7  (h]r8  (h]r9  (h]r:  (h	h�e]r;  (hh�e]r<  (hhe]r=  (h]r>  (h	h�e]r?  (hh�e]r@  (hhe]rA  (j�  ]rB  (h	h�e]rC  (hh�eeee]rD  (hhee]rE  (h!]rF  (h#h$e]rG  (h	j�  e]rH  (hh�e]rI  (h)heeej7  j7  j7  j7  j7  j7  ]rJ  (h]rK  (h]rL  (h]rM  (h	h�e]rN  (hh�e]rO  (hhe]rP  (h]rQ  (h	h�e]rR  (hh�e]rS  (hhe]rT  (j�  ]rU  (h	h�e]rV  (hh�eeee]rW  (hhee]rX  (h!]rY  (h#h$e]rZ  (h	j�  e]r[  (hh�e]r\  (h)heeejJ  jJ  jJ  jJ  jJ  jJ  ]r]  (h]r^  (h]r_  (h]r`  (h	h�e]ra  (hh�e]rb  (hhe]rc  (h]rd  (h	h�e]re  (hh�e]rf  (hhe]rg  (j�  ]rh  (h	h�e]ri  (hh�eeee]rj  (hhee]rk  (h!]rl  (h#h$e]rm  (h	j�  e]rn  (hh�e]ro  (h)heeej]  j]  j]  j]  j]  ]rp  (h]rq  (h]rr  (h]rs  (h	h�e]rt  (hh�e]ru  (hhe]rv  (h]rw  (h	h�e]rx  (hh�e]ry  (hhe]rz  (j�  ]r{  (h	h�e]r|  (hh�eeee]r}  (hhee]r~  (h!]r  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeejp  jp  jp  jp  jp  jp  jp  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r   (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej�  ]r  (h]r	  (h]r
  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej  j  j  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r   (hhe]r!  (h]r"  (h	h�e]r#  (hh�e]r$  (hhe]r%  (j�  ]r&  (h	h�e]r'  (hh�eeee]r(  (hhee]r)  (h!]r*  (h#h$e]r+  (h	j�  e]r,  (hh�e]r-  (h)heeej  j  j  j  j  j  j  j  j  j  ]r.  (h]r/  (h]r0  (h]r1  (h	h�e]r2  (hh�e]r3  (hhe]r4  (h]r5  (h	h�e]r6  (hh�e]r7  (hhe]r8  (j�  ]r9  (h	h�e]r:  (hh�eeee]r;  (hhee]r<  (h!]r=  (h#h$e]r>  (h	j�  e]r?  (hh�e]r@  (h)heeej.  j.  j.  ]rA  (h]rB  (h]rC  (h]rD  (h	h�e]rE  (hh�e]rF  (hhe]rG  (h]rH  (h	h�e]rI  (hh�e]rJ  (hhe]rK  (j�  ]rL  (h	h�e]rM  (hh�eeee]rN  (hhee]rO  (h!]rP  (h#h$e]rQ  (h	j�  e]rR  (hh�e]rS  (h)heeejA  jA  ]rT  (h]rU  (h]rV  (h]rW  (h	h�e]rX  (hh�e]rY  (hhe]rZ  (h]r[  (h	h�e]r\  (hh�e]r]  (hhe]r^  (j�  ]r_  (h	h�e]r`  (hh�eeee]ra  (hhee]rb  (h!]rc  (h#h$e]rd  (h	j�  e]re  (hh�e]rf  (h)heeejT  jT  ]rg  (h]rh  (h]ri  (h]rj  (h	h�e]rk  (hh�e]rl  (hhe]rm  (h]rn  (h	h�e]ro  (hh�e]rp  (hhe]rq  (j�  ]rr  (h	h�e]rs  (hh�eeee]rt  (hhee]ru  (h!]rv  (h#h$e]rw  (h	j�  e]rx  (hh�e]ry  (h)heeejg  jg  ]rz  (h]r{  (h]r|  (h]r}  (h	h�e]r~  (hh�e]r  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeejz  jz  jz  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r   (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r	  (j�  ]r
  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	j�  e]r  (hh�e]r  (h)heeej�  ]r  (h]r  (h]r  (h]r  (h	h�e]r  (hh�e]r  (hhe]r  (h]r  (h	he]r  (hh�e]r  (hhe]r  (j�  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r   (h!]r!  (h#h$e]r"  (h	j�  e]r#  (hh�e]r$  (h)heeej  j  j  j  ]r%  (h]r&  (h]r'  (h]r(  (h	h�e]r)  (hh�e]r*  (hhe]r+  (h]r,  (h	he]r-  (hh�e]r.  (hhe]r/  (j�  ]r0  (h	h�e]r1  (hh�eeee]r2  (hhee]r3  (h!]r4  (h#h$e]r5  (h	j�  e]r6  (hh�e]r7  (h)heeej%  ]r8  (h]r9  (h]r:  (h]r;  (h	h�e]r<  (hh�e]r=  (hhe]r>  (h]r?  (h	he]r@  (hh�e]rA  (hhe]rB  (j�  ]rC  (h	h�e]rD  (hh�eeee]rE  (hhee]rF  (h!]rG  (h#h$e]rH  (h	j�  e]rI  (hh�e]rJ  (h)heeej8  j8  ]rK  (h]rL  (h]rM  (h]rN  (h	h�e]rO  (hh�e]rP  (hhe]rQ  (h]rR  (h	he]rS  (hh�e]rT  (hhe]rU  (j�  ]rV  (h	h�e]rW  (hh�eeee]rX  (hhee]rY  (h!]rZ  (h#h$e]r[  (h	j�  e]r\  (hh�e]r]  (h)heee]r^  (h]r_  (h]r`  (h]ra  (h	h�e]rb  (hh�e]rc  (hhe]rd  (h]re  (h	he]rf  (hh�e]rg  (hhe]rh  (j�  ]ri  (h	h�e]rj  (hh�eeee]rk  (hhee]rl  (h!]rm  (h#h$e]rn  (h	j�  e]ro  (hh�e]rp  (h)heeej^  j^  ]rq  (h]rr  (h]rs  (h]rt  (h	h�e]ru  (hh�e]rv  (hhe]rw  (h]rx  (h	he]ry  (hh�e]rz  (hhe]r{  (j�  ]r|  (h	h�e]r}  (hh�eeee]r~  (hhee]r  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeejq  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (h]r�  (h]r�  (h]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (h]r�  (h	he]r�  (hh�e]r�  (hhe]r    (j�  ]r   (h	h�e]r   (hh�eeee]r   (hhee]r   (h!]r   (h#h$e]r   (h	j�  e]r   (hh�e]r   (h)heeej�  j�  j�  j�  j�  j�  j�  ]r	   (h]r
   (h]r   (h]r   (h	h�e]r   (hh�e]r   (hhe]r   (h]r   (h	he]r   (hh�e]r   (hhe]r   (j�  ]r   (h	h�e]r   (hh�eeee]r   (hhee]r   (h!]r   (h#h$e]r   (h	j�  e]r   (hh�e]r   (h)heee]r   (h]r   (h]r   (h]r   (h	h�e]r    (hh�e]r!   (hhe]r"   (h]r#   (h	he]r$   (hh�e]r%   (hhe]r&   (j�  ]r'   (h	h�e]r(   (hh�eeee]r)   (hhee]r*   (h!]r+   (h#h$e]r,   (h	j�  e]r-   (hh�e]r.   (h)heeej   j   j   j   j   j   j   ]r/   (h]r0   (h]r1   (h]r2   (h	h�e]r3   (hh�e]r4   (hhe]r5   (h]r6   (h	he]r7   (hh�e]r8   (hhe]r9   (j�  ]r:   (h	h�e]r;   (hh�eeee]r<   (hhee]r=   (h!]r>   (h#h$e]r?   (h	j�  e]r@   (hh�e]rA   (h)heeej/   j/   j/   j/   j/   ]rB   (h]rC   (h]rD   (h]rE   (h	h�e]rF   (hh�e]rG   (hhe]rH   (h]rI   (h	he]rJ   (hh�e]rK   (hhe]rL   (j�  ]rM   (h	h�e]rN   (hh�eeee]rO   (hhee]rP   (h!]rQ   (h#h$e]rR   (h	j�  e]rS   (hh�e]rT   (h)heeejB   ]rU   (h]rV   (h]rW   (h]rX   (h	h�e]rY   (hh�e]rZ   (hhe]r[   (h]r\   (h	he]r]   (hh�e]r^   (hhe]r_   (j�  ]r`   (h	h�e]ra   (hh�eeee]rb   (hhee]rc   (h!]rd   (h#h$e]re   (h	j�  e]rf   (hh�e]rg   (h)heeejU   ]rh   (h]ri   (h]rj   (h]rk   (h	h�e]rl   (hh�e]rm   (hhe]rn   (h]ro   (h	he]rp   (hh�e]rq   (hhe]rr   (j�  ]rs   (h	h�e]rt   (hh�eeee]ru   (hhee]rv   (h!]rw   (h#h$e]rx   (h	j�  e]ry   (hh�e]rz   (h)heeejh   jh   jh   jh   jh   ]r{   (h]r|   (h]r}   (h]r~   (h	h�e]r   (hh�e]r�   (hhe]r�   (h]r�   (h	he]r�   (hh�e]r�   (hhe]r�   (j�  ]r�   (h	h�e]r�   (hh�eeee]r�   (hhee]r�   (h!]r�   (h#h$e]r�   (h	j�  e]r�   (hh�e]r�   (h)heeej{   j{   ]r�   (h]r�   (h]r�   (h]r�   (h	h�e]r�   (hh�e]r�   (hhe]r�   (h]r�   (h	he]r�   (hh�e]r�   (hhe]r�   (j�  ]r�   (h	h�e]r�   (hh�eeee]r�   (hhee]r�   (h!]r�   (h#h$e]r�   (h	j�  e]r�   (hh�e]r�   (h)heeej�   j�   ]r�   (h]r�   (h]r�   (h]r�   (h	h�e]r�   (hh�e]r�   (hhe]r�   (h]r�   (h	he]r�   (hh�e]r�   (hhe]r�   (j�  ]r�   (h	h�e]r�   (hh�eeee]r�   (hhee]r�   (h!]r�   (h#h$e]r�   (h	j�  e]r�   (hh�e]r�   (h)heeej�   j�   ]r�   (h]r�   (h]r�   (h]r�   (h	h�e]r�   (hh�e]r�   (hhe]r�   (h]r�   (h	he]r�   (hh�e]r�   (hhe]r�   (j�  ]r�   (h	h�e]r�   (hh�eeee]r�   (hhee]r�   (h!]r�   (h#h$e]r�   (h	j�  e]r�   (hh�e]r�   (h)heee]r�   (h]r�   (h]r�   (h]r�   (h	h�e]r�   (hh�e]r�   (hhe]r�   (h]r�   (h	he]r�   (hh�e]r�   (hhe]r�   (j�  ]r�   (h	h�e]r�   (hh�eeee]r�   (hhee]r�   (h!]r�   (h#h$e]r�   (h	j�  e]r�   (hh�e]r�   (h)heeej�   j�   j�   ]r�   (h]r�   (h]r�   (h]r�   (h	h�e]r�   (hh�e]r�   (hhe]r�   (h]r�   (h	he]r�   (hh�e]r�   (hhe]r�   (j�  ]r�   (h	h�e]r�   (hh�eeee]r�   (hhee]r�   (h!]r�   (h#h$e]r�   (h	j�  e]r�   (hh�e]r�   (h)heeej�   j�   j�   j�   j�   j�   j�   j�   ]r�   (h]r�   (h]r�   (h]r�   (h	h�e]r�   (hh�e]r�   (hhe]r�   (h]r�   (h	he]r�   (hh�e]r�   (hhe]r�   (j�  ]r�   (h	h�e]r�   (hh�eeee]r�   (hhee]r�   (h!]r�   (h#h$e]r�   (h	j�  e]r�   (hh�e]r�   (h)heeej�   j�   j�   j�   ]r !  (h]r!  (h]r!  (h]r!  (h	h�e]r!  (hh�e]r!  (hhe]r!  (h]r!  (h	he]r!  (hh�e]r	!  (hhe]r
!  (j�  ]r!  (h	h�e]r!  (hh�eeee]r!  (hhee]r!  (h!]r!  (h#h$e]r!  (h	j�  e]r!  (hh�e]r!  (h)heeej !  j !  j !  ]r!  (h]r!  (h]r!  (h]r!  (h	h�e]r!  (hh�e]r!  (hhe]r!  (h]r!  (h	he]r!  (hh�e]r!  (hhe]r!  (j�  ]r!  (h	h�e]r!  (hh�eeee]r !  (hhee]r!!  (h!]r"!  (h#h$e]r#!  (h	j�  e]r$!  (hh�e]r%!  (h)heeej!  j!  j!  ]r&!  (h]r'!  (h]r(!  (h]r)!  (h	h�e]r*!  (hh�e]r+!  (hhe]r,!  (h]r-!  (h	he]r.!  (hh�e]r/!  (hhe]r0!  (j�  ]r1!  (h	h�e]r2!  (hh�eeee]r3!  (hhee]r4!  (h!]r5!  (h#h$e]r6!  (h	j�  e]r7!  (hh�e]r8!  (h)heeej&!  j&!  j&!  j&!  j&!  ]r9!  (h]r:!  (h]r;!  (h]r<!  (h	h�e]r=!  (hh�e]r>!  (hhe]r?!  (h]r@!  (h	he]rA!  (hh�e]rB!  (hhe]rC!  (j�  ]rD!  (h	h�e]rE!  (hh�eeee]rF!  (hhee]rG!  (h!]rH!  (h#h$e]rI!  (h	j�  e]rJ!  (hh�e]rK!  (h)heeej9!  j9!  j9!  ]rL!  (h]rM!  (h]rN!  (h]rO!  (h	h�e]rP!  (hh�e]rQ!  (hhe]rR!  (h]rS!  (h	he]rT!  (hh�e]rU!  (hhe]rV!  (j�  ]rW!  (h	h�e]rX!  (hh�eeee]rY!  (hhee]rZ!  (h!]r[!  (h#h$e]r\!  (h	j�  e]r]!  (hh�e]r^!  (h)heeejL!  jL!  jL!  jL!  jL!  ]r_!  (h]r`!  (h]ra!  (h]rb!  (h	h�e]rc!  (hh�e]rd!  (hhe]re!  (h]rf!  (h	he]rg!  (hh�e]rh!  (hhe]ri!  (X	   Next-Moverj!  ]rk!  (h	h�e]rl!  (hh�eeee]rm!  (hhee]rn!  (h!]ro!  (h#h$e]rp!  (h	j�  e]rq!  (hh�e]rr!  (h)heeej_!  j_!  ]rs!  (h]rt!  (h]ru!  (h]rv!  (h	h�e]rw!  (hh�e]rx!  (hhe]ry!  (h]rz!  (h	he]r{!  (hh�e]r|!  (hhe]r}!  (jj!  ]r~!  (h	h�e]r!  (hh�eeee]r�!  (hhee]r�!  (h!]r�!  (h#h$e]r�!  (h	j�  e]r�!  (hh�e]r�!  (h)heeejs!  js!  js!  js!  ]r�!  (h]r�!  (h]r�!  (h]r�!  (h	h�e]r�!  (hh�e]r�!  (hhe]r�!  (h]r�!  (h	he]r�!  (hh�e]r�!  (hhe]r�!  (jj!  ]r�!  (h	h�e]r�!  (hh�eeee]r�!  (hhee]r�!  (h!]r�!  (h#h$e]r�!  (h	j�  e]r�!  (hh�e]r�!  (h)heee]r�!  (h]r�!  (h]r�!  (h]r�!  (h	h�e]r�!  (hh�e]r�!  (hhe]r�!  (h]r�!  (h	he]r�!  (hh�e]r�!  (hhe]r�!  (jj!  ]r�!  (h	h�e]r�!  (hh�eeee]r�!  (hhee]r�!  (h!]r�!  (h#h$e]r�!  (h	j�  e]r�!  (hh�e]r�!  (h)heeej�!  ]r�!  (h]r�!  (h]r�!  (h]r�!  (h	h�e]r�!  (hh�e]r�!  (hhe]r�!  (h]r�!  (h	he]r�!  (hh�e]r�!  (hhe]r�!  (jj!  ]r�!  (h	h�e]r�!  (hh�eeee]r�!  (hhee]r�!  (h!]r�!  (h#h$e]r�!  (h	j�  e]r�!  (hh�e]r�!  (h)heeej�!  j�!  j�!  ]r�!  (h]r�!  (h]r�!  (h]r�!  (h	h�e]r�!  (hh�e]r�!  (hhe]r�!  (h]r�!  (h	he]r�!  (hh�e]r�!  (hhe]r�!  (jj!  ]r�!  (h	h�e]r�!  (hh�eeee]r�!  (hhee]r�!  (h!]r�!  (h#h$e]r�!  (h	j�  e]r�!  (hh�e]r�!  (h)heeej�!  j�!  j�!  j�!  ]r�!  (h]r�!  (h]r�!  (h]r�!  (h	h�e]r�!  (hh�e]r�!  (hhe]r�!  (h]r�!  (h	he]r�!  (hh�e]r�!  (hhe]r�!  (jj!  ]r�!  (h	h�e]r�!  (hh�eeee]r�!  (hhee]r�!  (h!]r�!  (h#h$e]r�!  (h	j�  e]r�!  (hh�e]r�!  (h)heeej�!  j�!  ]r�!  (h]r�!  (h]r�!  (h]r�!  (h	h�e]r�!  (hh�e]r�!  (hhe]r�!  (h]r�!  (h	he]r�!  (hh�e]r�!  (hhe]r�!  (jj!  ]r�!  (h	h�e]r�!  (hh�eeee]r�!  (hhee]r�!  (h!]r�!  (h#h$e]r�!  (h	j�  e]r�!  (hh�e]r�!  (h)heeej�!  j�!  j�!  j�!  ]r�!  (h]r�!  (h]r�!  (h]r�!  (h	h�e]r�!  (hh�e]r�!  (hhe]r�!  (h]r�!  (h	he]r "  (hh�e]r"  (hhe]r"  (jj!  ]r"  (h	h�e]r"  (hh�eeee]r"  (hhee]r"  (h!]r"  (h#h$e]r"  (h	j�  e]r	"  (hh�e]r
"  (h)heeej�!  ]r"  (h]r"  (h]r"  (h]r"  (h	h�e]r"  (hh�e]r"  (hhe]r"  (h]r"  (h	he]r"  (hh�e]r"  (hhe]r"  (jj!  ]r"  (h	h�e]r"  (hh�eeee]r"  (hhee]r"  (h!]r"  (h#h$e]r"  (h	j�  e]r"  (hh�e]r"  (h)heee]r"  (h]r"  (h]r "  (h]r!"  (h	h�e]r""  (hh�e]r#"  (hhe]r$"  (h]r%"  (h	he]r&"  (hh�e]r'"  (hhe]r("  (jj!  ]r)"  (h	h�e]r*"  (hh�eeee]r+"  (hhee]r,"  (h!]r-"  (h#h$e]r."  (h	j�  e]r/"  (hh�e]r0"  (h)heeej"  j"  ]r1"  (h]r2"  (h]r3"  (h]r4"  (h	h�e]r5"  (hh�e]r6"  (hhe]r7"  (h]r8"  (h	he]r9"  (hh�e]r:"  (hhe]r;"  (jj!  ]r<"  (h	h�e]r="  (hh�eeee]r>"  (hhee]r?"  (h!]r@"  (h#h$e]rA"  (h	j�  e]rB"  (hh�e]rC"  (h)heeej1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  j1"  ]rD"  (h]rE"  (h]rF"  (h]rG"  (h	h�e]rH"  (hh�e]rI"  (hhe]rJ"  (h]rK"  (h	he]rL"  (hh�e]rM"  (hhe]rN"  (jj!  ]rO"  (h	h�e]rP"  (hh�eeee]rQ"  (hhee]rR"  (h!]rS"  (h#h$e]rT"  (h	j�  e]rU"  (hh�e]rV"  (h)heeejD"  jD"  ]rW"  (h]rX"  (h]rY"  (h]rZ"  (h	h�e]r["  (hh�e]r\"  (hhe]r]"  (h]r^"  (h	he]r_"  (hh�e]r`"  (hhe]ra"  (jj!  ]rb"  (h	h�e]rc"  (hh�eeee]rd"  (hhee]re"  (h!]rf"  (h#h$e]rg"  (h	j�  e]rh"  (hh�e]ri"  (h)heeejW"  jW"  ]rj"  (h]rk"  (h]rl"  (h]rm"  (h	h�e]rn"  (hh�e]ro"  (hhe]rp"  (h]rq"  (h	he]rr"  (hh�e]rs"  (hhe]rt"  (jj!  ]ru"  (h	h�e]rv"  (hh�eeee]rw"  (hhee]rx"  (h!]ry"  (h#h$e]rz"  (h	j�  e]r{"  (hh�e]r|"  (h)heee]r}"  (h]r~"  (h]r"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (h]r�"  (h	he]r�"  (hh�e]r�"  (hhe]r�"  (jj!  ]r�"  (h	h�e]r�"  (hh�eeee]r�"  (hhee]r�"  (h!]r�"  (h#h$e]r�"  (h	j�  e]r�"  (hh�e]r�"  (h)heeej}"  j}"  j}"  j}"  ]r�"  (h]r�"  (h]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (jj!  ]r�"  (h	h�e]r�"  (hh�eeee]r�"  (hhee]r�"  (h!]r�"  (h#h$e]r�"  (h	j�  e]r�"  (hh�e]r�"  (h)heeej�"  j�"  j�"  j�"  j�"  j�"  j�"  ]r�"  (h]r�"  (h]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (jj!  ]r�"  (h	h�e]r�"  (hh�eeee]r�"  (hhee]r�"  (h!]r�"  (h#h$e]r�"  (h	j�  e]r�"  (hh�e]r�"  (h)heee]r�"  (h]r�"  (h]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (jj!  ]r�"  (h	h�e]r�"  (hh�eeee]r�"  (hhee]r�"  (h!]r�"  (h#h$e]r�"  (h	j�  e]r�"  (hh�e]r�"  (h)heeej�"  j�"  ]r�"  (h]r�"  (h]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (jj!  ]r�"  (h	h�e]r�"  (hh�eeee]r�"  (hhee]r�"  (h!]r�"  (h#h$e]r�"  (h	j�  e]r�"  (hh�e]r�"  (h)heeej�"  j�"  j�"  j�"  j�"  j�"  ]r�"  (h]r�"  (h]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (jj!  ]r�"  (h	h�e]r�"  (hh�eeee]r�"  (hhee]r�"  (h!]r�"  (h#h$e]r�"  (h	j�  e]r�"  (hh�e]r�"  (h)heeej�"  j�"  ]r�"  (h]r�"  (h]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (h]r�"  (h	h�e]r�"  (hh�e]r�"  (hhe]r�"  (jj!  ]r�"  (h	h�e]r�"  (hh�eeee]r�"  (hhee]r�"  (h!]r�"  (h#h$e]r�"  (h	j�  e]r #  (hh�e]r#  (h)heeej�"  j�"  j�"  j�"  ]r#  (h]r#  (h]r#  (h]r#  (h	h�e]r#  (hh�e]r#  (hhe]r#  (h]r	#  (h	h�e]r
#  (hh�e]r#  (hhe]r#  (jj!  ]r#  (h	h�e]r#  (hh�eeee]r#  (hhee]r#  (h!]r#  (h#h$e]r#  (h	j�  e]r#  (hh�e]r#  (h)heeej#  j#  j#  j#  j#  j#  j#  j#  j#  ]r#  (h]r#  (h]r#  (h]r#  (h	h�e]r#  (hh�e]r#  (hhe]r#  (h]r#  (h	h�e]r#  (hh�e]r#  (hhe]r#  (jj!  ]r #  (h	h�e]r!#  (hh�eeee]r"#  (hhee]r##  (h!]r$#  (h#h$e]r%#  (h	j�  e]r&#  (hh�e]r'#  (h)heeej#  j#  j#  j#  j#  j#  j#  ]r(#  (h]r)#  (h]r*#  (h]r+#  (h	h�e]r,#  (hh�e]r-#  (hhe]r.#  (h]r/#  (h	h�e]r0#  (hh�e]r1#  (hhe]r2#  (jj!  ]r3#  (h	h�e]r4#  (hh�eeee]r5#  (hhee]r6#  (h!]r7#  (h#h$e]r8#  (h	j�  e]r9#  (hh�e]r:#  (h)heee]r;#  (h]r<#  (h]r=#  (h]r>#  (h	h�e]r?#  (hh�e]r@#  (hhe]rA#  (h]rB#  (h	h�e]rC#  (hh�e]rD#  (hhe]rE#  (jj!  ]rF#  (h	h�e]rG#  (hh�eeee]rH#  (hhee]rI#  (h!]rJ#  (h#h$e]rK#  (h	j�  e]rL#  (hh�e]rM#  (h)heeej;#  j;#  j;#  j;#  j;#  j;#  j;#  j;#  j;#  ]rN#  (h]rO#  (h]rP#  (h]rQ#  (h	h�e]rR#  (hh�e]rS#  (hhe]rT#  (h]rU#  (h	h�e]rV#  (hh�e]rW#  (hhe]rX#  (jj!  ]rY#  (h	h�e]rZ#  (hh�eeee]r[#  (hhee]r\#  (h!]r]#  (h#h$e]r^#  (h	j�  e]r_#  (hh�e]r`#  (h)heeejN#  jN#  jN#  jN#  ]ra#  (h]rb#  (h]rc#  (h]rd#  (h	h�e]re#  (hh�e]rf#  (hhe]rg#  (h]rh#  (h	h�e]ri#  (hh�e]rj#  (hhe]rk#  (jj!  ]rl#  (h	h�e]rm#  (hh�eeee]rn#  (hhee]ro#  (h!]rp#  (h#h$e]rq#  (h	j�  e]rr#  (hh�e]rs#  (h)heeeja#  ja#  ja#  ja#  ]rt#  (h]ru#  (h]rv#  (h]rw#  (h	h�e]rx#  (hh�e]ry#  (hhe]rz#  (h]r{#  (h	h�e]r|#  (hh�e]r}#  (hhe]r~#  (jj!  ]r#  (h	h�e]r�#  (hh�eeee]r�#  (hhee]r�#  (h!]r�#  (h#h$e]r�#  (h	j�  e]r�#  (hh�e]r�#  (h)heeejt#  jt#  jt#  ]r�#  (h]r�#  (h]r�#  (h]r�#  (h	h�e]r�#  (hh�e]r�#  (hhe]r�#  (h]r�#  (h	h�e]r�#  (hh�e]r�#  (hhe]r�#  (jj!  ]r�#  (h	h�e]r�#  (hh�eeee]r�#  (hhee]r�#  (h!]r�#  (h#h$e]r�#  (h	j�  e]r�#  (hh�e]r�#  (h)heeej�#  ]r�#  (h]r�#  (h]r�#  (h]r�#  (h	h�e]r�#  (hh�e]r�#  (hhe]r�#  (h]r�#  (h	h�e]r�#  (hh�e]r�#  (hhe]r�#  (jj!  ]r�#  (h	h�e]r�#  (hh�eeee]r�#  (hhee]r�#  (h!]r�#  (h#h$e]r�#  (h	j�  e]r�#  (hh�e]r�#  (h)heeej�#  j�#  j�#  ]r�#  (h]r�#  (h]r�#  (h]r�#  (h	h�e]r�#  (hh�e]r�#  (hhe]r�#  (h]r�#  (h	h�e]r�#  (hh�e]r�#  (hhe]r�#  (jj!  ]r�#  (h	h�e]r�#  (hh�eeee]r�#  (hhee]r�#  (h!]r�#  (h#h$e]r�#  (h	j�  e]r�#  (hh�e]r�#  (h)heee]r�#  (h]r�#  (h]r�#  (h]r�#  (h	h�e]r�#  (hh�e]r�#  (hhe]r�#  (h]r�#  (h	h�e]r�#  (hh�e]r�#  (hhe]r�#  (jj!  ]r�#  (h	h�e]r�#  (hh�eeee]r�#  (hhee]r�#  (h!]r�#  (h#h$e]r�#  (h	j�  e]r�#  (hh�e]r�#  (h)heeej�#  j�#  ]r�#  (h]r�#  (h]r�#  (h]r�#  (h	h�e]r�#  (hh�e]r�#  (hhe]r�#  (h]r�#  (h	he]r�#  (hh�e]r�#  (hhe]r�#  (jj!  ]r�#  (h	h�e]r�#  (hh�eeee]r�#  (hhee]r�#  (h!]r�#  (h#h$e]r�#  (h	j�  e]r�#  (hh�e]r�#  (h)heeej�#  j�#  j�#  j�#  j�#  j�#  j�#  j�#  j�#  ]r�#  (h]r�#  (h]r�#  (h]r�#  (h	h�e]r�#  (hh�e]r�#  (hhe]r�#  (h]r�#  (h	he]r�#  (hh�e]r�#  (hhe]r�#  (jj!  ]r�#  (h	h�e]r�#  (hh�eeee]r�#  (hhee]r�#  (h!]r�#  (h#h$e]r�#  (h	j�  e]r�#  (hh�e]r�#  (h)heee]r�#  (h]r�#  (h]r�#  (h]r�#  (h	h�e]r�#  (hh�e]r�#  (hhe]r�#  (h]r $  (h	he]r$  (hh�e]r$  (hhe]r$  (jj!  ]r$  (h	h�e]r$  (hh�eeee]r$  (hhee]r$  (h!]r$  (h#h$e]r	$  (h	j�  e]r
$  (hh�e]r$  (h)heeej�#  j�#  j�#  j�#  j�#  ]r$  (h]r$  (h]r$  (h]r$  (h	h�e]r$  (hh�e]r$  (hhe]r$  (h]r$  (h	he]r$  (hh�e]r$  (hhe]r$  (jj!  ]r$  (h	h�e]r$  (hh�eeee]r$  (hhee]r$  (h!]r$  (h#h$e]r$  (h	j�  e]r$  (hh�e]r$  (h)heeej$  j$  ]r$  (h]r $  (h]r!$  (h]r"$  (h	h�e]r#$  (hh�e]r$$  (hhe]r%$  (h]r&$  (h	he]r'$  (hh�e]r($  (hhe]r)$  (jj!  ]r*$  (h	h�e]r+$  (hh�eeee]r,$  (hhee]r-$  (h!]r.$  (h#h$e]r/$  (h	j�  e]r0$  (hh�e]r1$  (h)heeej$  j$  j$  ]r2$  (h]r3$  (h]r4$  (h]r5$  (h	h�e]r6$  (hh�e]r7$  (hhe]r8$  (h]r9$  (h	he]r:$  (hh�e]r;$  (hhe]r<$  (jj!  ]r=$  (h	h�e]r>$  (hh�eeee]r?$  (hhee]r@$  (h!]rA$  (h#h$e]rB$  (h	j�  e]rC$  (hh�e]rD$  (h)heeej2$  j2$  j2$  ]rE$  (h]rF$  (h]rG$  (h]rH$  (h	h�e]rI$  (hh�e]rJ$  (hhe]rK$  (h]rL$  (h	he]rM$  (hh�e]rN$  (hhe]rO$  (jj!  ]rP$  (h	h�e]rQ$  (hh�eeee]rR$  (hhee]rS$  (h!]rT$  (h#h$e]rU$  (h	j�  e]rV$  (hh�e]rW$  (h)heeejE$  jE$  jE$  ]rX$  (h]rY$  (h]rZ$  (h]r[$  (h	h�e]r\$  (hh�e]r]$  (hhe]r^$  (h]r_$  (h	he]r`$  (hh�e]ra$  (hhe]rb$  (jj!  ]rc$  (h	h�e]rd$  (hh�eeee]re$  (hhee]rf$  (h!]rg$  (h#h$e]rh$  (h	j�  e]ri$  (hh�e]rj$  (h)heeejX$  jX$  jX$  jX$  ]rk$  (h]rl$  (h]rm$  (h]rn$  (h	h�e]ro$  (hh�e]rp$  (hhe]rq$  (h]rr$  (h	he]rs$  (hh�e]rt$  (hhe]ru$  (jj!  ]rv$  (h	h�e]rw$  (hh�eeee]rx$  (hhee]ry$  (h!]rz$  (h#h$e]r{$  (h	j�  e]r|$  (hh�e]r}$  (h)heeejk$  jk$  ]r~$  (h]r$  (h]r�$  (h]r�$  (h	h�e]r�$  (hh�e]r�$  (hhe]r�$  (h]r�$  (h	he]r�$  (hh�e]r�$  (hhe]r�$  (jj!  ]r�$  (h	h�e]r�$  (hh�eeee]r�$  (hhee]r�$  (h!]r�$  (h#h$e]r�$  (h	j�  e]r�$  (hh�e]r�$  (h)heeej~$  j~$  j~$  ]r�$  (h]r�$  (h]r�$  (h]r�$  (h	h�e]r�$  (hh�e]r�$  (hhe]r�$  (h]r�$  (h	he]r�$  (hh�e]r�$  (hhe]r�$  (jj!  ]r�$  (h	h�e]r�$  (hh�eeee]r�$  (hhee]r�$  (h!]r�$  (h#h$e]r�$  (h	j�  e]r�$  (hh�e]r�$  (h)heee]r�$  (h]r�$  (h]r�$  (h]r�$  (h	h�e]r�$  (hh�e]r�$  (hhe]r�$  (h]r�$  (h	he]r�$  (hh�e]r�$  (hhe]r�$  (jj!  ]r�$  (h	h�e]r�$  (hh�eeee]r�$  (hhee]r�$  (h!]r�$  (h#h$e]r�$  (h	j�  e]r�$  (hh�e]r�$  (h)heee]r�$  (h]r�$  (h]r�$  (h]r�$  (h	h�e]r�$  (hh�e]r�$  (hhe]r�$  (h]r�$  (h	he]r�$  (hh�e]r�$  (hhe]r�$  (jj!  ]r�$  (h	h�e]r�$  (hh�eeee]r�$  (hhee]r�$  (h!]r�$  (h#h$e]r�$  (h	j�  e]r�$  (hh�e]r�$  (h)heeej�$  j�$  j�$  ]r�$  (h]r�$  (h]r�$  (h]r�$  (h	h�e]r�$  (hh�e]r�$  (hhe]r�$  (h]r�$  (h	h�e]r�$  (hh�e]r�$  (hhe]r�$  (jj!  ]r�$  (h	h�e]r�$  (hh�eeee]r�$  (hhee]r�$  (h!]r�$  (h#h$e]r�$  (h	j�  e]r�$  (hh�e]r�$  (h)heee]r�$  (h]r�$  (h]r�$  (h]r�$  (h	h�e]r�$  (hh�e]r�$  (hhe]r�$  (h]r�$  (h	h�e]r�$  (hh�e]r�$  (hhe]r�$  (jj!  ]r�$  (h	h�e]r�$  (hh�eeee]r�$  (hhee]r�$  (h!]r�$  (h#h$e]r�$  (h	j�  e]r�$  (hh�e]r�$  (h)heee]r�$  (h]r�$  (h]r�$  (h]r�$  (h	h�e]r�$  (hh�e]r�$  (hhe]r�$  (h]r�$  (h	h�e]r�$  (hh�e]r�$  (hhe]r�$  (jj!  ]r�$  (h	h�e]r�$  (hh�eeee]r�$  (hhee]r�$  (h!]r�$  (h#h$e]r %  (h	j�  e]r%  (hh�e]r%  (h)heeej�$  j�$  j�$  j�$  j�$  j�$  j�$  ]r%  (h]r%  (h]r%  (h]r%  (h	h�e]r%  (hh�e]r%  (hhe]r	%  (h]r
%  (h	h�e]r%  (hh�e]r%  (hhe]r%  (jj!  ]r%  (h	h�e]r%  (hh�eeee]r%  (hhee]r%  (h!]r%  (h#h$e]r%  (h	j�  e]r%  (hh�e]r%  (h)heeej%  j%  j%  j%  j%  ]r%  (h]r%  (h]r%  (h]r%  (h	h�e]r%  (hh�e]r%  (hhe]r%  (h]r%  (h	h�e]r%  (hh�e]r%  (hhe]r %  (jj!  ]r!%  (h	h�e]r"%  (hh�eeee]r#%  (hhee]r$%  (h!]r%%  (h#h$e]r&%  (h	j�  e]r'%  (hh�e]r(%  (h)heeej%  j%  j%  ]r)%  (h]r*%  (h]r+%  (h]r,%  (h	h�e]r-%  (hh�e]r.%  (hhe]r/%  (h]r0%  (h	h�e]r1%  (hh�e]r2%  (hhe]r3%  (jj!  ]r4%  (h	h�e]r5%  (hh�eeee]r6%  (hhee]r7%  (h!]r8%  (h#h$e]r9%  (h	j�  e]r:%  (hh�e]r;%  (h)heeej)%  j)%  j)%  ]r<%  (h]r=%  (h]r>%  (h]r?%  (h	h�e]r@%  (hh�e]rA%  (hhe]rB%  (h]rC%  (h	h�e]rD%  (hh�e]rE%  (hhe]rF%  (jj!  ]rG%  (h	h�e]rH%  (hh�eeee]rI%  (hhee]rJ%  (h!]rK%  (h#h$e]rL%  (h	j�  e]rM%  (hh�e]rN%  (h)heeej<%  j<%  j<%  j<%  j<%  j<%  ]rO%  (h]rP%  (h]rQ%  (h]rR%  (h	h�e]rS%  (hh�e]rT%  (hhe]rU%  (h]rV%  (h	he]rW%  (hh�e]rX%  (hhe]rY%  (jj!  ]rZ%  (h	h�e]r[%  (hh�eeee]r\%  (hhee]r]%  (h!]r^%  (h#h$e]r_%  (h	j�  e]r`%  (hh�e]ra%  (h)heee]rb%  (h]rc%  (h]rd%  (h]re%  (h	h�e]rf%  (hh�e]rg%  (hhe]rh%  (h]ri%  (h	he]rj%  (hh�e]rk%  (hhe]rl%  (jj!  ]rm%  (h	h�e]rn%  (hh�eeee]ro%  (hhee]rp%  (h!]rq%  (h#h$e]rr%  (h	j�  e]rs%  (hh�e]rt%  (h)heeejb%  jb%  jb%  ]ru%  (h]rv%  (h]rw%  (h]rx%  (h	h�e]ry%  (hh�e]rz%  (hhe]r{%  (h]r|%  (h	he]r}%  (hh�e]r~%  (hhe]r%  (jj!  ]r�%  (h	h�e]r�%  (hh�eeee]r�%  (hhee]r�%  (h!]r�%  (h#h$e]r�%  (h	j�  e]r�%  (hh�e]r�%  (h)heeeju%  ju%  ju%  ju%  ju%  ]r�%  (h]r�%  (h]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (jj!  ]r�%  (h	h�e]r�%  (hh�eeee]r�%  (hhee]r�%  (h!]r�%  (h#h$e]r�%  (h	j�  e]r�%  (hh�e]r�%  (h)heee]r�%  (h]r�%  (h]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (jj!  ]r�%  (h	h�e]r�%  (hh�eeee]r�%  (hhee]r�%  (h!]r�%  (h#h$e]r�%  (h	j�  e]r�%  (hh�e]r�%  (h)heeej�%  j�%  j�%  j�%  ]r�%  (h]r�%  (h]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (jj!  ]r�%  (h	h�e]r�%  (hh�eeee]r�%  (hhee]r�%  (h!]r�%  (h#h$e]r�%  (h	j�  e]r�%  (hh�e]r�%  (h)heeej�%  j�%  j�%  ]r�%  (h]r�%  (h]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (jj!  ]r�%  (h	h�e]r�%  (hh�eeee]r�%  (hhee]r�%  (h!]r�%  (h#h$e]r�%  (h	j�  e]r�%  (hh�e]r�%  (h)heee]r�%  (h]r�%  (h]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (jj!  ]r�%  (h	h�e]r�%  (hh�eeee]r�%  (hhee]r�%  (h!]r�%  (h#h$e]r�%  (h	j�  e]r�%  (hh�e]r�%  (h)heee]r�%  (h]r�%  (h]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r�%  (jj!  ]r�%  (h	h�e]r�%  (hh�eeee]r�%  (hhee]r�%  (h!]r�%  (h#h$e]r�%  (h	j�  e]r�%  (hh�e]r�%  (h)heeej�%  ]r�%  (h]r�%  (h]r�%  (h]r�%  (h	h�e]r�%  (hh�e]r�%  (hhe]r &  (h]r&  (h	h�e]r&  (hh�e]r&  (hhe]r&  (jj!  ]r&  (h	h�e]r&  (hh�eeee]r&  (hhee]r&  (h!]r	&  (h#h$e]r
&  (h	j�  e]r&  (hh�e]r&  (h)heeej�%  j�%  j�%  j�%  j�%  ]r&  (h]r&  (h]r&  (h]r&  (h	h�e]r&  (hh�e]r&  (hhe]r&  (h]r&  (h	h�e]r&  (hh�e]r&  (hhe]r&  (jj!  ]r&  (h	h�e]r&  (hh�eeee]r&  (hhee]r&  (h!]r&  (h#h$e]r&  (h	j�  e]r&  (hh�e]r&  (h)heeej&  ]r &  (h]r!&  (h]r"&  (h]r#&  (h	h�e]r$&  (hh�e]r%&  (hhe]r&&  (h]r'&  (h	h�e]r(&  (hh�e]r)&  (hhe]r*&  (jj!  ]r+&  (h	h�e]r,&  (hh�eeee]r-&  (hhee]r.&  (h!]r/&  (h#h$e]r0&  (h	j�  e]r1&  (hh�e]r2&  (h)heeej &  j &  j &  j &  ]r3&  (h]r4&  (h]r5&  (h]r6&  (h	h�e]r7&  (hh�e]r8&  (hhe]r9&  (h]r:&  (h	h�e]r;&  (hh�e]r<&  (hhe]r=&  (jj!  ]r>&  (h	h�e]r?&  (hh�eeee]r@&  (hhee]rA&  (h!]rB&  (h#h$e]rC&  (h	j�  e]rD&  (hh�e]rE&  (h)heee]rF&  (h]rG&  (h]rH&  (h]rI&  (h	h�e]rJ&  (hh�e]rK&  (hhe]rL&  (h]rM&  (h	h�e]rN&  (hh�e]rO&  (hhe]rP&  (jj!  ]rQ&  (h	h�e]rR&  (hh�eeee]rS&  (hhee]rT&  (h!]rU&  (h#h$e]rV&  (h	j�  e]rW&  (hh�e]rX&  (h)heee]rY&  (h]rZ&  (h]r[&  (h]r\&  (h	h�e]r]&  (hh�e]r^&  (hhe]r_&  (h]r`&  (h	h�e]ra&  (hh�e]rb&  (hhe]rc&  (jj!  ]rd&  (h	h�e]re&  (hh�eeee]rf&  (hhee]rg&  (h!]rh&  (h#h$e]ri&  (h	j�  e]rj&  (hh�e]rk&  (h)heee]rl&  (h]rm&  (h]rn&  (h]ro&  (h	h�e]rp&  (hh�e]rq&  (hhe]rr&  (h]rs&  (h	h�e]rt&  (hh�e]ru&  (hhe]rv&  (jj!  ]rw&  (h	h�e]rx&  (hh�eeee]ry&  (hhee]rz&  (h!]r{&  (h#h$e]r|&  (h	j�  e]r}&  (hh�e]r~&  (h)heeejl&  jl&  jl&  jl&  jl&  ]r&  (h]r�&  (h]r�&  (h]r�&  (h	h�e]r�&  (hh�e]r�&  (hhe]r�&  (h]r�&  (h	h�e]r�&  (hh�e]r�&  (hhe]r�&  (jj!  ]r�&  (h	h�e]r�&  (hh�eeee]r�&  (hhee]r�&  (h!]r�&  (h#h$e]r�&  (h	j�  e]r�&  (hh�e]r�&  (h)heeej&  ]r�&  (h]r�&  (h]r�&  (h]r�&  (h	h�e]r�&  (hh�e]r�&  (hhe]r�&  (h]r�&  (h	h�e]r�&  (hh�e]r�&  (hhe]r�&  (jj!  ]r�&  (h	h�e]r�&  (hh�eeee]r�&  (hhee]r�&  (h!]r�&  (h#h$e]r�&  (h	j�  e]r�&  (hh�e]r�&  (h)heeej�&  ]r�&  (h]r�&  (h]r�&  (h]r�&  (h	h�e]r�&  (hh�e]r�&  (hhe]r�&  (h]r�&  (h	h�e]r�&  (hh�e]r�&  (hhe]r�&  (jj!  ]r�&  (h	h�e]r�&  (hh�eeee]r�&  (hhee]r�&  (h!]r�&  (h#h$e]r�&  (h	j�  e]r�&  (hh�e]r�&  (h)heeej�&  j�&  j�&  j�&  j�&  j�&  ]r�&  (h]r�&  (h]r�&  (h]r�&  (h	h�e]r�&  (hh�e]r�&  (hhe]r�&  (h]r�&  (h	h�e]r�&  (hh�e]r�&  (hhe]r�&  (jj!  ]r�&  (h	h�e]r�&  (hh�eeee]r�&  (hhee]r�&  (h!]r�&  (h#h$e]r�&  (h	j�  e]r�&  (hh�e]r�&  (h)heeej�&  ]r�&  (h]r�&  (h]r�&  (h]r�&  (h	h�e]r�&  (hh�e]r�&  (hhe]r�&  (h]r�&  (h	he]r�&  (hh�e]r�&  (hhe]r�&  (jj!  ]r�&  (h	h�e]r�&  (hh�eeee]r�&  (hhee]r�&  (h!]r�&  (h#h$e]r�&  (h	j�  e]r�&  (hh�e]r�&  (h)heeej�&  j�&  ]r�&  (h]r�&  (h]r�&  (h]r�&  (h	h�e]r�&  (hh�e]r�&  (hhe]r�&  (h]r�&  (h	he]r�&  (hh�e]r�&  (hhe]r�&  (jj!  ]r�&  (h	h�e]r�&  (hh�eeee]r�&  (hhee]r�&  (h!]r�&  (h#h$e]r�&  (h	j�  e]r�&  (hh�e]r�&  (h)heeej�&  ]r�&  (h]r�&  (h]r�&  (h]r�&  (h	h�e]r�&  (hh�e]r�&  (hhe]r�&  (h]r�&  (h	he]r�&  (hh�e]r�&  (hhe]r�&  (jj!  ]r�&  (h	h�e]r�&  (hh�eeee]r�&  (hhee]r�&  (h!]r '  (h#h$e]r'  (h	j�  e]r'  (hh�e]r'  (h)heeej�&  j�&  j�&  j�&  j�&  j�&  j�&  j�&  ]r'  (h]r'  (h]r'  (h]r'  (h	h�e]r'  (hh�e]r	'  (hhe]r
'  (h]r'  (h	he]r'  (hh�e]r'  (hhe]r'  (jj!  ]r'  (h	h�e]r'  (hh�eeee]r'  (hhee]r'  (h!]r'  (h#h$e]r'  (h	j�  e]r'  (hh�e]r'  (h)heeej'  ]r'  (h]r'  (h]r'  (h]r'  (h	h�e]r'  (hh�e]r'  (hhe]r'  (h]r'  (h	he]r'  (hh�e]r '  (hhe]r!'  (jj!  ]r"'  (h	h�e]r#'  (hh�eeee]r$'  (hhee]r%'  (h!]r&'  (h#h$e]r''  (h	j�  e]r('  (hh�e]r)'  (h)heeej'  j'  j'  j'  ]r*'  (h]r+'  (h]r,'  (h]r-'  (h	h�e]r.'  (hh�e]r/'  (hhe]r0'  (h]r1'  (h	he]r2'  (hh�e]r3'  (hhe]r4'  (jj!  ]r5'  (h	h�e]r6'  (hh�eeee]r7'  (hhee]r8'  (h!]r9'  (h#h$e]r:'  (h	j�  e]r;'  (hh�e]r<'  (h)heeej*'  j*'  ]r='  (h]r>'  (h]r?'  (h]r@'  (h	h�e]rA'  (hh�e]rB'  (hhe]rC'  (h]rD'  (h	he]rE'  (hh�e]rF'  (hhe]rG'  (jj!  ]rH'  (h	h�e]rI'  (hh�eeee]rJ'  (hhee]rK'  (h!]rL'  (h#h$e]rM'  (h	j�  e]rN'  (hh�e]rO'  (h)heeej='  j='  ]rP'  (h]rQ'  (h]rR'  (h]rS'  (h	h�e]rT'  (hh�e]rU'  (hhe]rV'  (h]rW'  (h	he]rX'  (hh�e]rY'  (hhe]rZ'  (jj!  ]r['  (h	h�e]r\'  (hh�eeee]r]'  (hhee]r^'  (h!]r_'  (h#h$e]r`'  (h	j�  e]ra'  (hh�e]rb'  (h)heeejP'  jP'  ]rc'  (h]rd'  (h]re'  (h]rf'  (h	h�e]rg'  (hh�e]rh'  (hhe]ri'  (h]rj'  (h	he]rk'  (hh�e]rl'  (hhe]rm'  (jj!  ]rn'  (h	h�e]ro'  (hh�eeee]rp'  (hhee]rq'  (h!]rr'  (h#h$e]rs'  (h	j�  e]rt'  (hh�e]ru'  (h)heeejc'  jc'  jc'  jc'  ]rv'  (h]rw'  (h]rx'  (h]ry'  (h	h�e]rz'  (hh�e]r{'  (hhe]r|'  (h]r}'  (h	he]r~'  (hh�e]r'  (hhe]r�'  (jj!  ]r�'  (h	h�e]r�'  (hh�eeee]r�'  (hhee]r�'  (h!]r�'  (h#h$e]r�'  (h	j�  e]r�'  (hh�e]r�'  (h)heeejv'  jv'  ]r�'  (h]r�'  (h]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r�'  (hhe]r�'  (h]r�'  (h	he]r�'  (hh�e]r�'  (hhe]r�'  (jj!  ]r�'  (h	h�e]r�'  (hh�eeee]r�'  (hhee]r�'  (h!]r�'  (h#h$e]r�'  (h	j�  e]r�'  (hh�e]r�'  (h)heeej�'  j�'  j�'  ]r�'  (h]r�'  (h]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r�'  (hhe]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r�'  (hhe]r�'  (jj!  ]r�'  (h	h�e]r�'  (hh�eeee]r�'  (hhee]r�'  (h!]r�'  (h#h$e]r�'  (h	j�  e]r�'  (hh�e]r�'  (h)heee]r�'  (h]r�'  (h]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r�'  (hhe]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r�'  (hhe]r�'  (jj!  ]r�'  (h	h�e]r�'  (hh�eeee]r�'  (hhee]r�'  (h!]r�'  (h#h$e]r�'  (h	j�  e]r�'  (hh�e]r�'  (h)heeej�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  j�'  ]r�'  (h]r�'  (h]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r�'  (hhe]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r�'  (hhe]r�'  (jj!  ]r�'  (h	h�e]r�'  (hh�eeee]r�'  (hhee]r�'  (h!]r�'  (h#h$e]r�'  (h	j�  e]r�'  (hh�e]r�'  (h)heeej�'  j�'  j�'  j�'  j�'  j�'  j�'  ]r�'  (h]r�'  (h]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r�'  (hhe]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r�'  (hhe]r�'  (jj!  ]r�'  (h	h�e]r�'  (hh�eeee]r�'  (hhee]r�'  (h!]r�'  (h#h$e]r�'  (h	j�  e]r�'  (hh�e]r�'  (h)heeej�'  j�'  ]r�'  (h]r�'  (h]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r�'  (hhe]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r�'  (hhe]r�'  (jj!  ]r�'  (h	h�e]r�'  (hh�eeee]r�'  (hhee]r�'  (h!]r�'  (h#h$e]r�'  (h	j�  e]r�'  (hh�e]r�'  (h)heeej�'  j�'  j�'  j�'  j�'  j�'  ]r�'  (h]r�'  (h]r�'  (h]r�'  (h	h�e]r�'  (hh�e]r (  (hhe]r(  (h]r(  (h	h�e]r(  (hh�e]r(  (hhe]r(  (jj!  ]r(  (h	h�e]r(  (hh�eeee]r(  (hhee]r	(  (h!]r
(  (h#h$e]r(  (h	j�  e]r(  (hh�e]r(  (h)heeej�'  j�'  ]r(  (h]r(  (h]r(  (h]r(  (h	h�e]r(  (hh�e]r(  (hhe]r(  (h]r(  (h	h�e]r(  (hh�e]r(  (hhe]r(  (jj!  ]r(  (h	h�e]r(  (hh�eeee]r(  (hhee]r(  (h!]r(  (h#h$e]r(  (h	j�  e]r(  (hh�e]r (  (h)heeej(  j(  j(  j(  j(  j(  j(  j(  j(  j(  j(  j(  j(  j(  j(  j(  j(  ]r!(  (h]r"(  (h]r#(  (h]r$(  (h	h�e]r%(  (hh�e]r&(  (hhe]r'(  (h]r((  (h	h�e]r)(  (hh�e]r*(  (hhe]r+(  (jj!  ]r,(  (h	h�e]r-(  (hh�eeee]r.(  (hhee]r/(  (h!]r0(  (h#h$e]r1(  (h	j�  e]r2(  (hh�e]r3(  (h)heeej!(  ]r4(  (h]r5(  (h]r6(  (h]r7(  (h	h�e]r8(  (hh�e]r9(  (hhe]r:(  (h]r;(  (h	h�e]r<(  (hh�e]r=(  (hhe]r>(  (jj!  ]r?(  (h	h�e]r@(  (hh�eeee]rA(  (hhee]rB(  (h!]rC(  (h#h$e]rD(  (h	j�  e]rE(  (hh�e]rF(  (h)heeej4(  j4(  j4(  j4(  ]rG(  (h]rH(  (h]rI(  (h]rJ(  (h	h�e]rK(  (hh�e]rL(  (hhe]rM(  (h]rN(  (h	h�e]rO(  (hh�e]rP(  (hhe]rQ(  (jj!  ]rR(  (h	h�e]rS(  (hh�eeee]rT(  (hhee]rU(  (h!]rV(  (h#h$e]rW(  (h	j�  e]rX(  (hh�e]rY(  (h)heeejG(  ]rZ(  (h]r[(  (h]r\(  (h]r](  (h	h�e]r^(  (hh�e]r_(  (hhe]r`(  (h]ra(  (h	h�e]rb(  (hh�e]rc(  (hhe]rd(  (jj!  ]re(  (h	h�e]rf(  (hh�eeee]rg(  (hhee]rh(  (h!]ri(  (h#h$e]rj(  (h	j�  e]rk(  (hh�e]rl(  (h)heeejZ(  jZ(  jZ(  ]rm(  (h]rn(  (h]ro(  (h]rp(  (h	h�e]rq(  (hh�e]rr(  (hhe]rs(  (h]rt(  (h	h�e]ru(  (hh�e]rv(  (hhe]rw(  (X	   Next-Moverx(  ]ry(  (h	h�e]rz(  (hh�eeee]r{(  (hhee]r|(  (h!]r}(  (h#h$e]r~(  (h	j�  e]r(  (hh�e]r�(  (h)heee]r�(  (h]r�(  (h]r�(  (h]r�(  (h	h�e]r�(  (hh�e]r�(  (hhe]r�(  (h]r�(  (h	he]r�(  (hh�e]r�(  (hhe]r�(  (jx(  ]r�(  (h	h�e]r�(  (hh�eeee]r�(  (hhee]r�(  (h!]r�(  (h#h$e]r�(  (h	j�  e]r�(  (hh�e]r�(  (h)heeej�(  ]r�(  (h]r�(  (h]r�(  (h]r�(  (h	h�e]r�(  (hh�e]r�(  (hhe]r�(  (h]r�(  (h	he]r�(  (hh�e]r�(  (hhe]r�(  (jx(  ]r�(  (h	h�e]r�(  (hh�eeee]r�(  (hhee]r�(  (h!]r�(  (h#h$e]r�(  (h	j�  e]r�(  (hh�e]r�(  (h)heeej�(  ]r�(  (h]r�(  (h]r�(  (h]r�(  (h	h�e]r�(  (hh�e]r�(  (hhe]r�(  (h]r�(  (h	he]r�(  (hh�e]r�(  (hhe]r�(  (jx(  ]r�(  (h	h�e]r�(  (hh�eeee]r�(  (hhee]r�(  (h!]r�(  (h#h$e]r�(  (h	j�  e]r�(  (hh�e]r�(  (h)heee]r�(  (h]r�(  (h]r�(  (h]r�(  (h	h�e]r�(  (hh�e]r�(  (hhe]r�(  (h]r�(  (h	he]r�(  (hh�e]r�(  (hhe]r�(  (jx(  ]r�(  (h	h�e]r�(  (hh�eeee]r�(  (hhee]r�(  (h!]r�(  (h#h$e]r�(  (h	j�  e]r�(  (hh�e]r�(  (h)heeej�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  j�(  ]r�(  (h]r�(  (h]r�(  (h]r�(  (h	h�e]r�(  (hh�e]r�(  (hhe]r�(  (h]r�(  (h	he]r�(  (hh�e]r�(  (hhe]r�(  (jx(  ]r�(  (h	h�e]r�(  (hh�eeee]r�(  (hhee]r�(  (h!]r�(  (h#h$e]r�(  (h	j�  e]r�(  (hh�e]r�(  (h)heee]r�(  (h]r�(  (h]r�(  (h]r�(  (h	h�e]r�(  (hh�e]r�(  (hhe]r�(  (h]r�(  (h	he]r�(  (hh�e]r�(  (hhe]r�(  (jx(  ]r�(  (h	h�e]r�(  (hh�eeee]r�(  (hhee]r�(  (h!]r�(  (h#h$e]r�(  (h	j�  e]r�(  (hh�e]r�(  (h)heeej�(  j�(  ]r�(  (h]r�(  (h]r�(  (h]r�(  (h	h�e]r�(  (hh�e]r�(  (hhe]r�(  (h]r�(  (h	he]r�(  (hh�e]r�(  (hhe]r�(  (jx(  ]r�(  (h	h�e]r�(  (hh�eeee]r )  (hhee]r)  (h!]r)  (h#h$e]r)  (h	j�  e]r)  (hh�e]r)  (h)heee]r)  (h]r)  (h]r)  (h]r	)  (h	h�e]r
)  (hh�e]r)  (hhe]r)  (h]r)  (h	he]r)  (hh�e]r)  (hhe]r)  (jx(  ]r)  (h	h�e]r)  (hh�eeee]r)  (hhee]r)  (h!]r)  (h#h$e]r)  (h	j�  e]r)  (hh�e]r)  (h)heeej)  j)  j)  ]r)  (h]r)  (h]r)  (h]r)  (h	h�e]r)  (hh�e]r)  (hhe]r)  (h]r )  (h	he]r!)  (hh�e]r")  (hhe]r#)  (jx(  ]r$)  (h	h�e]r%)  (hh�eeee]r&)  (hhee]r')  (h!]r()  (h#h$e]r))  (h	j�  e]r*)  (hh�e]r+)  (h)heeej)  j)  j)  j)  ]r,)  (h]r-)  (h]r.)  (h]r/)  (h	h�e]r0)  (hh�e]r1)  (hhe]r2)  (h]r3)  (h	he]r4)  (hh�e]r5)  (hhe]r6)  (jx(  ]r7)  (h	h�e]r8)  (hh�eeee]r9)  (hhee]r:)  (h!]r;)  (h#h$e]r<)  (h	j�  e]r=)  (hh�e]r>)  (h)heeej,)  j,)  j,)  j,)  j,)  j,)  j,)  j,)  j,)  ]r?)  (h]r@)  (h]rA)  (h]rB)  (h	h�e]rC)  (hh�e]rD)  (hhe]rE)  (h]rF)  (h	he]rG)  (hh�e]rH)  (hhe]rI)  (jx(  ]rJ)  (h	h�e]rK)  (hh�eeee]rL)  (hhee]rM)  (h!]rN)  (h#h$e]rO)  (h	j�  e]rP)  (hh�e]rQ)  (h)heeej?)  j?)  j?)  j?)  ]rR)  (h]rS)  (h]rT)  (h]rU)  (h	h�e]rV)  (hh�e]rW)  (hhe]rX)  (h]rY)  (h	he]rZ)  (hh�e]r[)  (hhe]r\)  (jx(  ]r])  (h	h�e]r^)  (hh�eeee]r_)  (hhee]r`)  (h!]ra)  (h#h$e]rb)  (h	j�  e]rc)  (hh�e]rd)  (h)heeejR)  jR)  jR)  ]re)  (h]rf)  (h]rg)  (h]rh)  (h	h�e]ri)  (hh�e]rj)  (hhe]rk)  (h]rl)  (h	he]rm)  (hh�e]rn)  (hhe]ro)  (jx(  ]rp)  (h	h�e]rq)  (hh�eeee]rr)  (hhee]rs)  (h!]rt)  (h#h$e]ru)  (h	j�  e]rv)  (hh�e]rw)  (h)heeeje)  je)  je)  ]rx)  (h]ry)  (h]rz)  (h]r{)  (h	h�e]r|)  (hh�e]r})  (hhe]r~)  (h]r)  (h	he]r�)  (hh�e]r�)  (hhe]r�)  (jx(  ]r�)  (h	h�e]r�)  (hh�eeee]r�)  (hhee]r�)  (h!]r�)  (h#h$e]r�)  (h	j�  e]r�)  (hh�e]r�)  (h)heeejx)  jx)  ]r�)  (h]r�)  (h]r�)  (h]r�)  (h	h�e]r�)  (hh�e]r�)  (hhe]r�)  (h]r�)  (h	he]r�)  (hh�e]r�)  (hhe]r�)  (jx(  ]r�)  (h	h�e]r�)  (hh�eeee]r�)  (hhee]r�)  (h!]r�)  (h#h$e]r�)  (h	j�  e]r�)  (hh�e]r�)  (h)heeej�)  j�)  j�)  j�)  j�)  j�)  j�)  ]r�)  (h]r�)  (h]r�)  (h]r�)  (h	h�e]r�)  (hh�e]r�)  (hhe]r�)  (h]r�)  (h	he]r�)  (hh�e]r�)  (hhe]r�)  (jx(  ]r�)  (h	h�e]r�)  (hh�eeee]r�)  (hhee]r�)  (h!]r�)  (h#h$e]r�)  (h	j�  e]r�)  (hh�e]r�)  (h)heeej�)  ]r�)  (h]r�)  (h]r�)  (h]r�)  (h	h�e]r�)  (hh�e]r�)  (hhe]r�)  (h]r�)  (h	he]r�)  (hh�e]r�)  (hhe]r�)  (jx(  ]r�)  (h	h�e]r�)  (hh�eeee]r�)  (hhee]r�)  (h!]r�)  (h#h$e]r�)  (h	j�  e]r�)  (hh�e]r�)  (h)heeej�)  j�)  j�)  ]r�)  (h]r�)  (h]r�)  (h]r�)  (h	h�e]r�)  (hh�e]r�)  (hhe]r�)  (h]r�)  (h	he]r�)  (hh�e]r�)  (hhe]r�)  (jx(  ]r�)  (h	h�e]r�)  (hh�eeee]r�)  (hhee]r�)  (h!]r�)  (h#h$e]r�)  (h	j�  e]r�)  (hh�e]r�)  (h)heeej�)  j�)  ]r�)  (h]r�)  (h]r�)  (h]r�)  (h	h�e]r�)  (hh�e]r�)  (hhe]r�)  (h]r�)  (h	he]r�)  (hh�e]r�)  (hhe]r�)  (jx(  ]r�)  (h	h�e]r�)  (hh�eeee]r�)  (hhee]r�)  (h!]r�)  (h#h$e]r�)  (h	j�  e]r�)  (hh�e]r�)  (h)heee]r�)  (h]r�)  (h]r�)  (h]r�)  (h	h�e]r�)  (hh�e]r�)  (hhe]r�)  (h]r�)  (h	he]r�)  (hh�e]r�)  (hhe]r�)  (jx(  ]r�)  (h	h�e]r�)  (hh�eeee]r�)  (hhee]r�)  (h!]r�)  (h#h$e]r�)  (h	j�  e]r�)  (hh�e]r�)  (h)heeej�)  j�)  ]r�)  (h]r�)  (h]r�)  (h]r *  (h	h�e]r*  (hh�e]r*  (hhe]r*  (h]r*  (h	he]r*  (hh�e]r*  (hhe]r*  (jx(  ]r*  (h	h�e]r	*  (hh�eeee]r
*  (hhee]r*  (h!]r*  (h#h$e]r*  (h	j�  e]r*  (hh�e]r*  (h)heeej�)  ]r*  (h]r*  (h]r*  (h]r*  (h	h�e]r*  (hh�e]r*  (hhe]r*  (h]r*  (h	he]r*  (hh�e]r*  (hhe]r*  (jx(  ]r*  (h	h�e]r*  (hh�eeee]r*  (hhee]r*  (h!]r*  (h#h$e]r *  (h	j�  e]r!*  (hh�e]r"*  (h)heeej*  ]r#*  (h]r$*  (h]r%*  (h]r&*  (h	h�e]r'*  (hh�e]r(*  (hhe]r)*  (h]r**  (h	he]r+*  (hh�e]r,*  (hhe]r-*  (jx(  ]r.*  (h	h�e]r/*  (hh�eeee]r0*  (hhee]r1*  (h!]r2*  (h#h$e]r3*  (h	j�  e]r4*  (hh�e]r5*  (h)heeej#*  ]r6*  (h]r7*  (h]r8*  (h]r9*  (h	h�e]r:*  (hh�e]r;*  (hhe]r<*  (h]r=*  (h	he]r>*  (hh�e]r?*  (hhe]r@*  (jx(  ]rA*  (h	h�e]rB*  (hh�eeee]rC*  (hhee]rD*  (h!]rE*  (h#h$e]rF*  (h	j�  e]rG*  (hh�e]rH*  (h)heee]rI*  (h]rJ*  (h]rK*  (h]rL*  (h	h�e]rM*  (hh�e]rN*  (hhe]rO*  (h]rP*  (h	he]rQ*  (hh�e]rR*  (hhe]rS*  (jx(  ]rT*  (h	h�e]rU*  (hh�eeee]rV*  (hhee]rW*  (h!]rX*  (h#h$e]rY*  (h	j�  e]rZ*  (hh�e]r[*  (h)heeejI*  jI*  jI*  jI*  jI*  jI*  ]r\*  (h]r]*  (h]r^*  (h]r_*  (h	h�e]r`*  (hh�e]ra*  (hhe]rb*  (h]rc*  (h	he]rd*  (hh�e]re*  (hhe]rf*  (jx(  ]rg*  (h	h�e]rh*  (hh�eeee]ri*  (hhee]rj*  (h!]rk*  (h#h$e]rl*  (h	j�  e]rm*  (hh�e]rn*  (h)heeej\*  j\*  ]ro*  (h]rp*  (h]rq*  (h]rr*  (h	h�e]rs*  (hh�e]rt*  (hhe]ru*  (h]rv*  (h	he]rw*  (hh�e]rx*  (hhe]ry*  (jx(  ]rz*  (h	h�e]r{*  (hh�eeee]r|*  (hhee]r}*  (h!]r~*  (h#h$e]r*  (h	j�  e]r�*  (hh�e]r�*  (h)heeejo*  jo*  jo*  jo*  ]r�*  (h]r�*  (h]r�*  (h]r�*  (h	h�e]r�*  (hh�e]r�*  (hhe]r�*  (h]r�*  (h	he]r�*  (hh�e]r�*  (hhe]r�*  (jx(  ]r�*  (h	h�e]r�*  (hh�eeee]r�*  (hhee]r�*  (h!]r�*  (h#h$e]r�*  (h	j�  e]r�*  (hh�e]r�*  (h)heee]r�*  (h]r�*  (h]r�*  (h]r�*  (h	h�e]r�*  (hh�e]r�*  (hhe]r�*  (h]r�*  (h	he]r�*  (hh�e]r�*  (hhe]r�*  (jx(  ]r�*  (h	h�e]r�*  (hh�eeee]r�*  (hhee]r�*  (h!]r�*  (h#h$e]r�*  (h	j�  e]r�*  (hh�e]r�*  (h)heeej�*  j�*  j�*  ]r�*  (h]r�*  (h]r�*  (h]r�*  (h	h�e]r�*  (hh�e]r�*  (hhe]r�*  (h]r�*  (h	he]r�*  (hh�e]r�*  (hhe]r�*  (jx(  ]r�*  (h	h�e]r�*  (hh�eeee]r�*  (hhee]r�*  (h!]r�*  (h#h$e]r�*  (h	j�  e]r�*  (hh�e]r�*  (h)heeej�*  j�*  ]r�*  (h]r�*  (h]r�*  (h]r�*  (h	h�e]r�*  (hh�e]r�*  (hhe]r�*  (h]r�*  (h	he]r�*  (hh�e]r�*  (hhe]r�*  (jx(  ]r�*  (h	h�e]r�*  (hh�eeee]r�*  (hhee]r�*  (h!]r�*  (h#h$e]r�*  (h	j�  e]r�*  (hh�e]r�*  (h)heeej�*  j�*  j�*  j�*  ]r�*  (h]r�*  (h]r�*  (h]r�*  (h	h�e]r�*  (hh�e]r�*  (hhe]r�*  (h]r�*  (h	he]r�*  (hh�e]r�*  (hhe]r�*  (jx(  ]r�*  (h	h�e]r�*  (hh�eeee]r�*  (hhee]r�*  (h!]r�*  (h#h$e]r�*  (h	j�  e]r�*  (hh�e]r�*  (h)heeej�*  j�*  j�*  j�*  ]r�*  (h]r�*  (h]r�*  (h]r�*  (h	h�e]r�*  (hh�e]r�*  (hhe]r�*  (h]r�*  (h	he]r�*  (hh�e]r�*  (hhe]r�*  (jx(  ]r�*  (h	h�e]r�*  (hh�eeee]r�*  (hhee]r�*  (h!]r�*  (h#h$e]r�*  (h	j�  e]r�*  (hh�e]r�*  (h)heeej�*  ]r�*  (h]r�*  (h]r�*  (h]r�*  (h	h�e]r�*  (hh�e]r�*  (hhe]r�*  (h]r�*  (h	he]r�*  (hh�e]r�*  (hhe]r�*  (jx(  ]r�*  (h	h�e]r +  (hh�eeee]r+  (hhee]r+  (h!]r+  (h#h$e]r+  (h	j�  e]r+  (hh�e]r+  (h)heeej�*  j�*  j�*  j�*  ]r+  (h]r+  (h]r	+  (h]r
+  (h	h�e]r+  (hh�e]r+  (hhe]r+  (h]r+  (h	he]r+  (hh�e]r+  (hhe]r+  (jx(  ]r+  (h	h�e]r+  (hh�eeee]r+  (hhee]r+  (h!]r+  (h#h$e]r+  (h	j�  e]r+  (hh�e]r+  (h)heee]r+  (h]r+  (h]r+  (h]r+  (h	h�e]r+  (hh�e]r+  (hhe]r +  (h]r!+  (h	he]r"+  (hh�e]r#+  (hhe]r$+  (jx(  ]r%+  (h	h�e]r&+  (hh�eeee]r'+  (hhee]r(+  (h!]r)+  (h#h$e]r*+  (h	j�  e]r++  (hh�e]r,+  (h)heeej+  j+  ]r-+  (h]r.+  (h]r/+  (h]r0+  (h	h�e]r1+  (hh�e]r2+  (hhe]r3+  (h]r4+  (h	he]r5+  (hh�e]r6+  (hhe]r7+  (jx(  ]r8+  (h	h�e]r9+  (hh�eeee]r:+  (hhee]r;+  (h!]r<+  (h#h$e]r=+  (h	j�  e]r>+  (hh�e]r?+  (h)heeej-+  j-+  j-+  j-+  j-+  j-+  j-+  j-+  j-+  ]r@+  (h]rA+  (h]rB+  (h]rC+  (h	h�e]rD+  (hh�e]rE+  (hhe]rF+  (h]rG+  (h	he]rH+  (hh�e]rI+  (hhe]rJ+  (jx(  ]rK+  (h	h�e]rL+  (hh�eeee]rM+  (hhee]rN+  (h!]rO+  (h#h$e]rP+  (h	j�  e]rQ+  (hh�e]rR+  (h)heeej@+  j@+  j@+  j@+  j@+  j@+  j@+  j@+  j@+  ]rS+  (h]rT+  (h]rU+  (h]rV+  (h	h�e]rW+  (hh�e]rX+  (hhe]rY+  (h]rZ+  (h	he]r[+  (hh�e]r\+  (hhe]r]+  (jx(  ]r^+  (h	h�e]r_+  (hh�eeee]r`+  (hhee]ra+  (h!]rb+  (h#h$e]rc+  (h	j�  e]rd+  (hh�e]re+  (h)heeejS+  jS+  jS+  jS+  ]rf+  (h]rg+  (h]rh+  (h]ri+  (h	h�e]rj+  (hh�e]rk+  (hhe]rl+  (h]rm+  (h	he]rn+  (hh�e]ro+  (hhe]rp+  (jx(  ]rq+  (h	h�e]rr+  (hh�eeee]rs+  (hhee]rt+  (h!]ru+  (h#h$e]rv+  (h	j�  e]rw+  (hh�e]rx+  (h)heeejf+  jf+  jf+  ]ry+  (h]rz+  (h]r{+  (h]r|+  (h	h�e]r}+  (hh�e]r~+  (hhe]r+  (h]r�+  (h	he]r�+  (hh�e]r�+  (hhe]r�+  (jx(  ]r�+  (h	h�e]r�+  (hh�eeee]r�+  (hhee]r�+  (h!]r�+  (h#h$e]r�+  (h	j�  e]r�+  (hh�e]r�+  (h)heeejy+  jy+  jy+  jy+  ]r�+  (h]r�+  (h]r�+  (h]r�+  (h	h�e]r�+  (hh�e]r�+  (hhe]r�+  (h]r�+  (h	he]r�+  (hh�e]r�+  (hhe]r�+  (jx(  ]r�+  (h	h�e]r�+  (hh�eeee]r�+  (hhee]r�+  (h!]r�+  (h#h$e]r�+  (h	j�  e]r�+  (hh�e]r�+  (h)heeej�+  j�+  j�+  ]r�+  (h]r�+  (h]r�+  (h]r�+  (h	h�e]r�+  (hh�e]r�+  (hhe]r�+  (h]r�+  (h	he]r�+  (hh�e]r�+  (hhe]r�+  (jx(  ]r�+  (h	h�e]r�+  (hh�eeee]r�+  (hhee]r�+  (h!]r�+  (h#h$e]r�+  (h	j�  e]r�+  (hh�e]r�+  (h)heeej�+  j�+  ]r�+  (h]r�+  (h]r�+  (h]r�+  (h	h�e]r�+  (hh�e]r�+  (hhe]r�+  (h]r�+  (h	he]r�+  (hh�e]r�+  (hhe]r�+  (jx(  ]r�+  (h	h�e]r�+  (hh�eeee]r�+  (hhee]r�+  (h!]r�+  (h#h$e]r�+  (h	j�  e]r�+  (hh�e]r�+  (h)heeej�+  j�+  j�+  ]r�+  (h]r�+  (h]r�+  (h]r�+  (h	h�e]r�+  (hh�e]r�+  (hhe]r�+  (h]r�+  (h	he]r�+  (hh�e]r�+  (hhe]r�+  (jx(  ]r�+  (h	h�e]r�+  (hh�eeee]r�+  (hhee]r�+  (h!]r�+  (h#h$e]r�+  (h	j�  e]r�+  (hh�e]r�+  (h)heeej�+  j�+  j�+  ]r�+  (h]r�+  (h]r�+  (h]r�+  (h	h�e]r�+  (hh�e]r�+  (hhe]r�+  (h]r�+  (h	he]r�+  (hh�e]r�+  (hhe]r�+  (jx(  ]r�+  (h	h�e]r�+  (hh�eeee]r�+  (hhee]r�+  (h!]r�+  (h#h$e]r�+  (h	j�  e]r�+  (hh�e]r�+  (h)heeej�+  j�+  j�+  ]r�+  (h]r�+  (h]r�+  (h]r�+  (h	h�e]r�+  (hh�e]r�+  (hhe]r�+  (h]r�+  (h	he]r�+  (hh�e]r�+  (hhe]r�+  (jx(  ]r�+  (h	h�e]r�+  (hh�eeee]r�+  (hhee]r�+  (h!]r�+  (h#h$e]r�+  (h	j�  e]r�+  (hh�e]r�+  (h)heeej�+  j�+  ]r�+  (h]r�+  (h]r ,  (h]r,  (h	h�e]r,  (hh�e]r,  (hhe]r,  (h]r,  (h	he]r,  (hh�e]r,  (hhe]r,  (jx(  ]r	,  (h	h�e]r
,  (hh�eeee]r,  (hhee]r,  (h!]r,  (h#h$e]r,  (h	j�  e]r,  (hh�e]r,  (h)heeej�+  ]r,  (h]r,  (h]r,  (h]r,  (h	h�e]r,  (hh�e]r,  (hhe]r,  (h]r,  (h	he]r,  (hh�e]r,  (hhe]r,  (jx(  ]r,  (h	h�e]r,  (hh�eeee]r,  (hhee]r,  (h!]r ,  (h#h$e]r!,  (h	j�  e]r",  (hh�e]r#,  (h)heee]r$,  (h]r%,  (h]r&,  (h]r',  (h	h�e]r(,  (hh�e]r),  (hhe]r*,  (h]r+,  (h	he]r,,  (hh�e]r-,  (hhe]r.,  (jx(  ]r/,  (h	h�e]r0,  (hh�eeee]r1,  (hhee]r2,  (h!]r3,  (h#h$e]r4,  (h	j�  e]r5,  (hh�e]r6,  (h)heeej$,  j$,  j$,  j$,  j$,  j$,  j$,  ]r7,  (h]r8,  (h]r9,  (h]r:,  (h	h�e]r;,  (hh�e]r<,  (hhe]r=,  (h]r>,  (h	h�e]r?,  (hh�e]r@,  (hhe]rA,  (jx(  ]rB,  (h	h�e]rC,  (hh�eeee]rD,  (hhee]rE,  (h!]rF,  (h#h$e]rG,  (h	j�  e]rH,  (hh�e]rI,  (h)heeej7,  ]rJ,  (h]rK,  (h]rL,  (h]rM,  (h	h�e]rN,  (hh�e]rO,  (hhe]rP,  (h]rQ,  (h	h�e]rR,  (hh�e]rS,  (hhe]rT,  (jx(  ]rU,  (h	h�e]rV,  (hh�eeee]rW,  (hhee]rX,  (h!]rY,  (h#h$e]rZ,  (h	j�  e]r[,  (hh�e]r\,  (h)heeejJ,  jJ,  jJ,  jJ,  jJ,  ]r],  (h]r^,  (h]r_,  (h]r`,  (h	h�e]ra,  (hh�e]rb,  (hhe]rc,  (h]rd,  (h	h�e]re,  (hh�e]rf,  (hhe]rg,  (jx(  ]rh,  (h	h�e]ri,  (hh�eeee]rj,  (hhee]rk,  (h!]rl,  (h#h$e]rm,  (h	j�  e]rn,  (hh�e]ro,  (h)heeej],  ]rp,  (h]rq,  (h]rr,  (h]rs,  (h	h�e]rt,  (hh�e]ru,  (hhe]rv,  (h]rw,  (h	h�e]rx,  (hh�e]ry,  (hhe]rz,  (jx(  ]r{,  (h	h�e]r|,  (hh�eeee]r},  (hhee]r~,  (h!]r,  (h#h$e]r�,  (h	j�  e]r�,  (hh�e]r�,  (h)heeejp,  jp,  ]r�,  (h]r�,  (h]r�,  (h]r�,  (h	h�e]r�,  (hh�e]r�,  (hhe]r�,  (h]r�,  (h	h�e]r�,  (hh�e]r�,  (hhe]r�,  (jx(  ]r�,  (h	h�e]r�,  (hh�eeee]r�,  (hhee]r�,  (h!]r�,  (h#h$e]r�,  (h	j�  e]r�,  (hh�e]r�,  (h)heeej�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  j�,  ]r�,  (h]r�,  (h]r�,  (h]r�,  (h	h�e]r�,  (hh�e]r�,  (hhe]r�,  (h]r�,  (h	h�e]r�,  (hh�e]r�,  (hhe]r�,  (jx(  ]r�,  (h	h�e]r�,  (hh�eeee]r�,  (hhee]r�,  (h!]r�,  (h#h$e]r�,  (h	j�  e]r�,  (hh�e]r�,  (h)heeee(]r�,  (h]r�,  (h]r�,  (h]r�,  (h	h�e]r�,  (hh�e]r�,  (hhe]r�,  (h]r�,  (h	he]r�,  (hh�e]r�,  (hhe]r�,  (jx(  ]r�,  (h	h�e]r�,  (hh�eeee]r�,  (hhee]r�,  (h!]r�,  (h#h$e]r�,  (h	j�  e]r�,  (hh�e]r�,  (h)heeee]r�,  (]r�,  (X   Normr�,  ]r�,  (X   Oblr�,  ]r�,  (X   Movedr�,  ]r�,  (h	j�  e]r�,  (hX   anyr�,  e]r�,  (hhe]r�,  (X   Movedr�,  ]r�,  (h	X   anyr�,  e]r�,  (hX   triangler�,  e]r�,  (hhe]r�,  (X	   Next-Mover�,  ]r�,  (h	he]r�,  (hX   squarer�,  eeee]r�,  (hheeej�,  j�,  ]r�,  (j�,  ]r�,  (j�,  ]r�,  (j�,  ]r�,  (h	j�  e]r�,  (hj�,  e]r�,  (hhe]r�,  (j�,  ]r�,  (h	j�,  e]r�,  (hj�,  e]r�,  (hhe]r�,  (j�,  ]r�,  (h	he]r�,  (hh�eeee]r�,  (hheeej�,  j�,  ]r�,  (j�,  ]r�,  (j�,  ]r�,  (j�,  ]r�,  (h	j�  e]r�,  (hj�,  e]r�,  (hhe]r�,  (j�,  ]r�,  (h	j�,  e]r�,  (hj�,  e]r�,  (hhe]r�,  (j�,  ]r�,  (h	he]r�,  (hh�eeee]r�,  (hheee]r�,  (j�,  ]r�,  (j�,  ]r�,  (j�,  ]r�,  (h	j�  e]r�,  (hj�,  e]r�,  (hhe]r�,  (j�,  ]r�,  (h	j�,  e]r�,  (hh�e]r�,  (hhe]r�,  (j�,  ]r�,  (h	he]r�,  (hh�eeee]r�,  (hheeej�,  ]r�,  (j�,  ]r�,  (j�,  ]r -  (j�,  ]r-  (h	j�  e]r-  (hj�,  e]r-  (hhe]r-  (j�,  ]r-  (h	j�,  e]r-  (hh�e]r-  (hhe]r-  (j�,  ]r	-  (h	he]r
-  (hh�eeee]r-  (hheee]r-  (j�,  ]r-  (j�,  ]r-  (j�,  ]r-  (h	j�  e]r-  (hh�e]r-  (hhe]r-  (j�,  ]r-  (h	j�,  e]r-  (hh�e]r-  (hhe]r-  (j�,  ]r-  (h	he]r-  (hh�eeee]r-  (hheeej-  ]r-  (j�,  ]r-  (j�,  ]r-  (j�,  ]r-  (h	j�  e]r-  (hh�e]r-  (hhe]r -  (j�,  ]r!-  (h	j�,  e]r"-  (hh�e]r#-  (hhe]r$-  (j�,  ]r%-  (h	h�e]r&-  (hh�eeee]r'-  (hheeej-  j-  j-  j-  j-  j-  ]r(-  (j�,  ]r)-  (j�,  ]r*-  (j�,  ]r+-  (h	j�  e]r,-  (hh�e]r--  (hhe]r.-  (j�,  ]r/-  (h	j�,  e]r0-  (hh�e]r1-  (hhe]r2-  (j�,  ]r3-  (h	h�e]r4-  (hh�eeee]r5-  (hheeej(-  ]r6-  (j�,  ]r7-  (j�,  ]r8-  (j�,  ]r9-  (h	j�  e]r:-  (hh�e]r;-  (hhe]r<-  (j�,  ]r=-  (h	j�,  e]r>-  (hh�e]r?-  (hhe]r@-  (j�,  ]rA-  (h	h�e]rB-  (hh�eeee]rC-  (hheeej6-  j6-  j6-  j6-  ]rD-  (j�,  ]rE-  (j�,  ]rF-  (j�,  ]rG-  (h	j�  e]rH-  (hh�e]rI-  (hhe]rJ-  (j�,  ]rK-  (h	j�,  e]rL-  (hh�e]rM-  (hhe]rN-  (j�,  ]rO-  (h	h�e]rP-  (hh�eeee]rQ-  (hheeejD-  jD-  ]rR-  (j�,  ]rS-  (j�,  ]rT-  (j�,  ]rU-  (h	j�  e]rV-  (hh�e]rW-  (hhe]rX-  (j�,  ]rY-  (h	j�,  e]rZ-  (hh�e]r[-  (hhe]r\-  (j�,  ]r]-  (h	h�e]r^-  (hh�eeee]r_-  (hheeejR-  ]r`-  (j�,  ]ra-  (j�,  ]rb-  (j�,  ]rc-  (h	j�  e]rd-  (hh�e]re-  (hhe]rf-  (j�,  ]rg-  (h	j�,  e]rh-  (hh�e]ri-  (hhe]rj-  (j�,  ]rk-  (h	h�e]rl-  (hh�eeee]rm-  (hheeej`-  j`-  j`-  ]rn-  (j�,  ]ro-  (j�,  ]rp-  (j�,  ]rq-  (h	j�  e]rr-  (hh�e]rs-  (hhe]rt-  (j�,  ]ru-  (h	j�,  e]rv-  (hh�e]rw-  (hhe]rx-  (j�,  ]ry-  (h	h�e]rz-  (hh�eeee]r{-  (hheee]r|-  (j�,  ]r}-  (j�,  ]r~-  (j�,  ]r-  (h	j�  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	j�,  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	h�e]r�-  (hh�eeee]r�-  (hheee]r�-  (j�,  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (h	j�  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	j�,  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	h�e]r�-  (hh�eeee]r�-  (hheeej�-  j�-  j�-  j�-  j�-  j�-  j�-  j�-  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (h	j�  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	j�,  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	h�e]r�-  (hh�eeee]r�-  (hheee]r�-  (j�,  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (h	j�  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	j�,  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	h�e]r�-  (hh�eeee]r�-  (hheee]r�-  (j�,  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (h	j�  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	j�,  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	h�e]r�-  (hh�eeee]r�-  (hheeej�-  j�-  j�-  j�-  j�-  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (h	j�  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	j�,  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	h�e]r�-  (hh�eeee]r�-  (hheeej�-  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (h	j�  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	j�,  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	h�e]r�-  (hh�eeee]r�-  (hheeej�-  j�-  j�-  j�-  j�-  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (h	j�  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	j�,  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	h�e]r�-  (hh�eeee]r�-  (hheeej�-  j�-  j�-  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (h	j�  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	j�,  e]r�-  (hh�e]r�-  (hhe]r�-  (j�,  ]r�-  (h	h�e]r�-  (hh�eeee]r�-  (hheeej�-  j�-  j�-  j�-  j�-  j�-  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (j�,  ]r�-  (h	j�  e]r�-  (hh�e]r�-  (hhe]r .  (j�,  ]r.  (h	j�,  e]r.  (hh�e]r.  (hhe]r.  (j�,  ]r.  (h	h�e]r.  (hh�eeee]r.  (hheeej�-  j�-  j�-  ]r.  (j�,  ]r	.  (j�,  ]r
.  (j�,  ]r.  (h	j�  e]r.  (hh�e]r.  (hhe]r.  (j�,  ]r.  (h	j�,  e]r.  (hh�e]r.  (hhe]r.  (j�,  ]r.  (h	h�e]r.  (hh�eeee]r.  (hheee]r.  (j�,  ]r.  (j�,  ]r.  (j�,  ]r.  (h	j�  e]r.  (hh�e]r.  (hhe]r.  (j�,  ]r.  (h	j�,  e]r.  (hh�e]r.  (hhe]r .  (X	   Next-Mover!.  ]r".  (h	h�e]r#.  (hh�eeee]r$.  (hheee]r%.  (j�,  ]r&.  (j�,  ]r'.  (j�,  ]r(.  (h	j�  e]r).  (hh�e]r*.  (hhe]r+.  (j�,  ]r,.  (h	j�,  e]r-.  (hh�e]r..  (hhe]r/.  (j!.  ]r0.  (h	he]r1.  (hh�eeee]r2.  (hheeej%.  j%.  j%.  j%.  ]r3.  (j�,  ]r4.  (j�,  ]r5.  (j�,  ]r6.  (h	j�  e]r7.  (hh�e]r8.  (hhe]r9.  (j�,  ]r:.  (h	j�,  e]r;.  (hh�e]r<.  (hhe]r=.  (j!.  ]r>.  (h	he]r?.  (hh�eeee]r@.  (hheeej3.  j3.  j3.  ]rA.  (j�,  ]rB.  (j�,  ]rC.  (j�,  ]rD.  (h	j�  e]rE.  (hh�e]rF.  (hhe]rG.  (j�,  ]rH.  (h	j�,  e]rI.  (hh�e]rJ.  (hhe]rK.  (j!.  ]rL.  (h	h�e]rM.  (hh�eeee]rN.  (hheee]rO.  (j�,  ]rP.  (j�,  ]rQ.  (j�,  ]rR.  (h	j�  e]rS.  (hh�e]rT.  (hhe]rU.  (j�,  ]rV.  (h	j�,  e]rW.  (hh�e]rX.  (hhe]rY.  (X	   Next-MoverZ.  ]r[.  (h	he]r\.  (hh�eeee]r].  (hheeejO.  jO.  jO.  ]r^.  (j�,  ]r_.  (j�,  ]r`.  (j�,  ]ra.  (h	j�  e]rb.  (hh�e]rc.  (hhe]rd.  (j�,  ]re.  (h	j�,  e]rf.  (hh�e]rg.  (hhe]rh.  (jZ.  ]ri.  (h	he]rj.  (hh�eeee]rk.  (hheeej^.  ]rl.  (j�,  ]rm.  (j�,  ]rn.  (j�,  ]ro.  (h	j�  e]rp.  (hh�e]rq.  (hhe]rr.  (j�,  ]rs.  (h	j�,  e]rt.  (hh�e]ru.  (hhe]rv.  (jZ.  ]rw.  (h	he]rx.  (hh�eeee]ry.  (hheeejl.  jl.  jl.  jl.  ]rz.  (j�,  ]r{.  (j�,  ]r|.  (j�,  ]r}.  (h	j�  e]r~.  (hh�e]r.  (hhe]r�.  (j�,  ]r�.  (h	j�,  e]r�.  (hh�e]r�.  (hhe]r�.  (jZ.  ]r�.  (h	h�e]r�.  (hh�eeee]r�.  (hheeejz.  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (h	j�  e]r�.  (hh�e]r�.  (hhe]r�.  (j�,  ]r�.  (h	j�,  e]r�.  (hh�e]r�.  (hhe]r�.  (jZ.  ]r�.  (h	h�e]r�.  (hh�eeee]r�.  (hheeej�.  j�.  j�.  j�.  j�.  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (h	j�  e]r�.  (hh�e]r�.  (hhe]r�.  (j�,  ]r�.  (h	j�,  e]r�.  (hh�e]r�.  (hhe]r�.  (jZ.  ]r�.  (h	h�e]r�.  (hh�eeee]r�.  (hheeej�.  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (h	j�  e]r�.  (hh�e]r�.  (hhe]r�.  (j�,  ]r�.  (h	j�,  e]r�.  (hh<e]r�.  (hhe]r�.  (jZ.  ]r�.  (h	h�e]r�.  (hh�eeee]r�.  (hheee]r�.  (j�,  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (h	j�  e]r�.  (hh�e]r�.  (hhe]r�.  (j�,  ]r�.  (h	j�,  e]r�.  (hh�e]r�.  (hhe]r�.  (jZ.  ]r�.  (h	h�e]r�.  (hh�eeee]r�.  (hheeej�.  j�.  j�.  j�.  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (h	j�  e]r�.  (hh�e]r�.  (hhe]r�.  (j�,  ]r�.  (h	j�,  e]r�.  (hh�e]r�.  (hhe]r�.  (jZ.  ]r�.  (h	h�e]r�.  (hh�eeee]r�.  (hheeej�.  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (h	j�  e]r�.  (hh�e]r�.  (hhe]r�.  (j�,  ]r�.  (h	j�,  e]r�.  (hh�e]r�.  (hhe]r�.  (jZ.  ]r�.  (h	h�e]r�.  (hh�eeee]r�.  (hheeej�.  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (h	j�  e]r�.  (hh�e]r�.  (hhe]r�.  (j�,  ]r�.  (h	j�,  e]r�.  (hh�e]r�.  (hhe]r�.  (jZ.  ]r�.  (h	h�e]r�.  (hh�eeee]r�.  (hheeej�.  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (h	j�  e]r�.  (hh�e]r�.  (hhe]r�.  (j�,  ]r�.  (h	j�,  e]r�.  (hh�e]r�.  (hhe]r�.  (jZ.  ]r�.  (h	h�e]r�.  (hh�eeee]r�.  (hheeej�.  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (j�,  ]r�.  (h	j�  e]r�.  (hh�e]r�.  (hhe]r�.  (j�,  ]r�.  (h	j�,  e]r /  (hh�e]r/  (hhe]r/  (jZ.  ]r/  (h	h�e]r/  (hh�eeee]r/  (hheeej�.  j�.  ]r/  (j�,  ]r/  (j�,  ]r/  (j�,  ]r	/  (h	j�  e]r
/  (hh�e]r/  (hhe]r/  (j�,  ]r/  (h	j�,  e]r/  (hh�e]r/  (hhe]r/  (jZ.  ]r/  (h	h�e]r/  (hh�eeee]r/  (hheee]r/  (j�,  ]r/  (j�,  ]r/  (j�,  ]r/  (h	j�  e]r/  (hh�e]r/  (hhe]r/  (j�,  ]r/  (h	j�,  e]r/  (hh�e]r/  (hhe]r/  (jZ.  ]r/  (h	h�e]r /  (hh�eeee]r!/  (hheeej/  j/  j/  j/  j/  ]r"/  (j�,  ]r#/  (j�,  ]r$/  (j�,  ]r%/  (h	j�  e]r&/  (hh�e]r'/  (hhe]r(/  (j�,  ]r)/  (h	j�,  e]r*/  (hh�e]r+/  (hhe]r,/  (jZ.  ]r-/  (h	h�e]r./  (hh�eeee]r//  (hheee]r0/  (j�,  ]r1/  (j�,  ]r2/  (j�,  ]r3/  (h	j�  e]r4/  (hh�e]r5/  (hhe]r6/  (j�,  ]r7/  (h	j�,  e]r8/  (hh�e]r9/  (hhe]r:/  (jZ.  ]r;/  (h	h�e]r</  (hh�eeee]r=/  (hheeej0/  ]r>/  (j�,  ]r?/  (j�,  ]r@/  (j�,  ]rA/  (h	j�  e]rB/  (hh�e]rC/  (hhe]rD/  (j�,  ]rE/  (h	j�,  e]rF/  (hh�e]rG/  (hhe]rH/  (jZ.  ]rI/  (h	h�e]rJ/  (hh�eeee]rK/  (hheee]rL/  (j�,  ]rM/  (j�,  ]rN/  (j�,  ]rO/  (h	j�  e]rP/  (hh�e]rQ/  (hhe]rR/  (j�,  ]rS/  (h	j�,  e]rT/  (hh�e]rU/  (hhe]rV/  (jZ.  ]rW/  (h	h�e]rX/  (hh�eeee]rY/  (hheeejL/  jL/  jL/  jL/  ]rZ/  (j�,  ]r[/  (j�,  ]r\/  (j�,  ]r]/  (h	j�  e]r^/  (hh�e]r_/  (hhe]r`/  (j�,  ]ra/  (h	h�e]rb/  (hh�e]rc/  (hhe]rd/  (jZ.  ]re/  (h	h�e]rf/  (hh�eeee]rg/  (hheeejZ/  jZ/  jZ/  ]rh/  (j�,  ]ri/  (j�,  ]rj/  (j�,  ]rk/  (h	j�  e]rl/  (hh�e]rm/  (hhe]rn/  (j�,  ]ro/  (h	h�e]rp/  (hh�e]rq/  (hhe]rr/  (jZ.  ]rs/  (h	h�e]rt/  (hh�eeee]ru/  (hheee]rv/  (j�,  ]rw/  (j�,  ]rx/  (j�,  ]ry/  (h	j�  e]rz/  (hh�e]r{/  (hhe]r|/  (j�,  ]r}/  (h	h�e]r~/  (hh�e]r/  (hhe]r�/  (jZ.  ]r�/  (h	h�e]r�/  (hh�eeee]r�/  (hheee]r�/  (j�,  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (h	j�  e]r�/  (hh�e]r�/  (hhe]r�/  (j�,  ]r�/  (h	h�e]r�/  (hh�e]r�/  (hhe]r�/  (jZ.  ]r�/  (h	h�e]r�/  (hh�eeee]r�/  (hheee]r�/  (j�,  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (h	j�  e]r�/  (hh�e]r�/  (hhe]r�/  (j�,  ]r�/  (h	h�e]r�/  (hh�e]r�/  (hhe]r�/  (jZ.  ]r�/  (h	h�e]r�/  (hh�eeee]r�/  (hheeej�/  j�/  j�/  j�/  j�/  j�/  j�/  j�/  j�/  j�/  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (h	j�  e]r�/  (hh�e]r�/  (hhe]r�/  (j�,  ]r�/  (h	h�e]r�/  (hh�e]r�/  (hhe]r�/  (jZ.  ]r�/  (h	he]r�/  (hh�eeee]r�/  (hheeej�/  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (h	j�  e]r�/  (hh�e]r�/  (hhe]r�/  (j�,  ]r�/  (h	h�e]r�/  (hh�e]r�/  (hhe]r�/  (jZ.  ]r�/  (h	he]r�/  (hh�eeee]r�/  (hheeej�/  j�/  j�/  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (h	j�  e]r�/  (hh�e]r�/  (hhe]r�/  (j�,  ]r�/  (h	h�e]r�/  (hh�e]r�/  (hhe]r�/  (jZ.  ]r�/  (h	h�e]r�/  (hh�eeee]r�/  (hheee]r�/  (j�,  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (h	j�  e]r�/  (hh�e]r�/  (hhe]r�/  (j�,  ]r�/  (h	h�e]r�/  (hh�e]r�/  (hhe]r�/  (jZ.  ]r�/  (h	h�e]r�/  (hh�eeee]r�/  (hheee]r�/  (j�,  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (h	j�  e]r�/  (hh�e]r�/  (hhe]r�/  (j�,  ]r�/  (h	h�e]r�/  (hh�e]r�/  (hhe]r�/  (jZ.  ]r�/  (h	h�e]r�/  (hh�eeee]r�/  (hheeej�/  j�/  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (h	j�  e]r�/  (hh�e]r�/  (hhe]r�/  (j�,  ]r�/  (h	h�e]r�/  (hh�e]r�/  (hhe]r�/  (jZ.  ]r�/  (h	h�e]r�/  (hh�eeee]r�/  (hheee]r�/  (j�,  ]r�/  (j�,  ]r�/  (j�,  ]r�/  (h	j�  e]r�/  (hh�e]r�/  (hhe]r�/  (j�,  ]r�/  (h	h�e]r�/  (hh�e]r�/  (hhe]r�/  (jZ.  ]r�/  (h	h�e]r 0  (hh�eeee]r0  (hheee]r0  (j�,  ]r0  (j�,  ]r0  (j�,  ]r0  (h	j�  e]r0  (hh�e]r0  (hhe]r0  (j�,  ]r	0  (h	h�e]r
0  (hh�e]r0  (hhe]r0  (jZ.  ]r0  (h	h�e]r0  (hh�eeee]r0  (hheee]r0  (j�,  ]r0  (j�,  ]r0  (j�,  ]r0  (h	j�  e]r0  (hh�e]r0  (hhe]r0  (j�,  ]r0  (h	h�e]r0  (hh�e]r0  (hhe]r0  (jZ.  ]r0  (h	h�e]r0  (hh�eeee]r0  (hheeej0  j0  j0  ]r0  (j�,  ]r0  (j�,  ]r 0  (j�,  ]r!0  (h	j�  e]r"0  (hh�e]r#0  (hhe]r$0  (j�,  ]r%0  (h	h�e]r&0  (hh�e]r'0  (hhe]r(0  (jZ.  ]r)0  (h	h�e]r*0  (hh�eeee]r+0  (hheeej0  ]r,0  (j�,  ]r-0  (j�,  ]r.0  (j�,  ]r/0  (h	j�  e]r00  (hh�e]r10  (hhe]r20  (j�,  ]r30  (h	h�e]r40  (hh�e]r50  (hhe]r60  (jZ.  ]r70  (h	h�e]r80  (hh�eeee]r90  (hheeej,0  j,0  j,0  ]r:0  (j�,  ]r;0  (j�,  ]r<0  (j�,  ]r=0  (h	j�  e]r>0  (hh�e]r?0  (hhe]r@0  (j�,  ]rA0  (h	h�e]rB0  (hh�e]rC0  (hhe]rD0  (jZ.  ]rE0  (h	h�e]rF0  (hh�eeee]rG0  (hheeej:0  j:0  j:0  j:0  j:0  ]rH0  (j�,  ]rI0  (j�,  ]rJ0  (j�,  ]rK0  (h	j�  e]rL0  (hh�e]rM0  (hhe]rN0  (j�,  ]rO0  (h	h�e]rP0  (hh�e]rQ0  (hhe]rR0  (jZ.  ]rS0  (h	h�e]rT0  (hh�eeee]rU0  (hheeejH0  ]rV0  (j�,  ]rW0  (j�,  ]rX0  (j�,  ]rY0  (h	j�  e]rZ0  (hh�e]r[0  (hhe]r\0  (j�,  ]r]0  (h	h�e]r^0  (hh�e]r_0  (hhe]r`0  (jZ.  ]ra0  (h	h�e]rb0  (hh�eeee]rc0  (hheee]rd0  (j�,  ]re0  (j�,  ]rf0  (j�,  ]rg0  (h	j�  e]rh0  (hh�e]ri0  (hhe]rj0  (j�,  ]rk0  (h	h�e]rl0  (hh�e]rm0  (hhe]rn0  (X	   Next-Movero0  ]rp0  (h	h�e]rq0  (hh�eeee]rr0  (hheee]rs0  (j�,  ]rt0  (j�,  ]ru0  (j�,  ]rv0  (h	j�  e]rw0  (hh�e]rx0  (hhe]ry0  (j�,  ]rz0  (h	h�e]r{0  (hh�e]r|0  (hhe]r}0  (X	   Next-Mover~0  ]r0  (h	he]r�0  (hh�eeee]r�0  (hheee]r�0  (j�,  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (h	j�  e]r�0  (hh�e]r�0  (hhe]r�0  (j�,  ]r�0  (h	h�e]r�0  (hh�e]r�0  (hhe]r�0  (j~0  ]r�0  (h	he]r�0  (hh�eeee]r�0  (hheee]r�0  (j�,  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (h	j�  e]r�0  (hh�e]r�0  (hhe]r�0  (j�,  ]r�0  (h	h�e]r�0  (hh�e]r�0  (hhe]r�0  (j~0  ]r�0  (h	he]r�0  (hh�eeee]r�0  (hheeej�0  j�0  j�0  j�0  j�0  j�0  j�0  j�0  j�0  j�0  j�0  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (h	j�  e]r�0  (hh�e]r�0  (hhe]r�0  (j�,  ]r�0  (h	h�e]r�0  (hh�e]r�0  (hhe]r�0  (j~0  ]r�0  (h	he]r�0  (hh�eeee]r�0  (hheeej�0  j�0  j�0  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (h	j�  e]r�0  (hh�e]r�0  (hhe]r�0  (j�,  ]r�0  (h	h�e]r�0  (hh�e]r�0  (hhe]r�0  (j~0  ]r�0  (h	he]r�0  (hh�eeee]r�0  (hheeej�0  j�0  j�0  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (h	j�  e]r�0  (hh�e]r�0  (hhe]r�0  (j�,  ]r�0  (h	h�e]r�0  (hh�e]r�0  (hhe]r�0  (j~0  ]r�0  (h	he]r�0  (hh�eeee]r�0  (hheee]r�0  (j�,  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (h	j�  e]r�0  (hh�e]r�0  (hhe]r�0  (j�,  ]r�0  (h	h�e]r�0  (hh�e]r�0  (hhe]r�0  (j~0  ]r�0  (h	he]r�0  (hh�eeee]r�0  (hheeej�0  j�0  j�0  j�0  j�0  j�0  j�0  j�0  j�0  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (h	j�  e]r�0  (hh�e]r�0  (hhe]r�0  (j�,  ]r�0  (h	h�e]r�0  (hh�e]r�0  (hhe]r�0  (j~0  ]r�0  (h	he]r�0  (hh�eeee]r�0  (hheeej�0  j�0  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (h	j�  e]r�0  (hh�e]r�0  (hhe]r�0  (j�,  ]r�0  (h	h�e]r�0  (hh�e]r�0  (hhe]r�0  (j~0  ]r�0  (h	he]r�0  (hh�eeee]r�0  (hheeej�0  j�0  j�0  j�0  j�0  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (j�,  ]r�0  (h	j�  e]r�0  (hh�e]r�0  (hhe]r�0  (j�,  ]r�0  (h	h�e]r�0  (hh�e]r�0  (hhe]r�0  (j~0  ]r�0  (h	he]r�0  (hh�eeee]r�0  (hheeej�0  j�0  j�0  j�0  j�0  j�0  j�0  j�0  j�0  ]r 1  (j�,  ]r1  (j�,  ]r1  (j�,  ]r1  (h	h�e]r1  (hh�e]r1  (hhe]r1  (j�,  ]r1  (h	h�e]r1  (hh�e]r	1  (hhe]r
1  (j~0  ]r1  (h	he]r1  (hh�eeee]r1  (hheeej 1  j 1  j 1  ]r1  (j�,  ]r1  (j�,  ]r1  (j�,  ]r1  (h	h�e]r1  (hh�e]r1  (hhe]r1  (j�,  ]r1  (h	h�e]r1  (hh�e]r1  (hhe]r1  (j~0  ]r1  (h	he]r1  (hh�eeee]r1  (hheeej1  j1  j1  j1  j1  j1  j1  ]r1  (j�,  ]r1  (j�,  ]r1  (j�,  ]r1  (h	h�e]r 1  (hh�e]r!1  (hhe]r"1  (j�,  ]r#1  (h	h�e]r$1  (hh�e]r%1  (hhe]r&1  (j~0  ]r'1  (h	he]r(1  (hh�eeee]r)1  (hheeej1  j1  ]r*1  (j�,  ]r+1  (j�,  ]r,1  (j�,  ]r-1  (h	h�e]r.1  (hh�e]r/1  (hhe]r01  (j�,  ]r11  (h	h�e]r21  (hh�e]r31  (hhe]r41  (j~0  ]r51  (h	he]r61  (hh�eeee]r71  (hheeej*1  j*1  j*1  j*1  j*1  j*1  ]r81  (j�,  ]r91  (j�,  ]r:1  (j�,  ]r;1  (h	h�e]r<1  (hh�e]r=1  (hhe]r>1  (j�,  ]r?1  (h	h�e]r@1  (hh�e]rA1  (hhe]rB1  (j~0  ]rC1  (h	he]rD1  (hh�eeee]rE1  (hheeej81  j81  ]rF1  (j�,  ]rG1  (j�,  ]rH1  (j�,  ]rI1  (h	j�  e]rJ1  (hh�e]rK1  (hhe]rL1  (j�,  ]rM1  (h	h�e]rN1  (hh�e]rO1  (hhe]rP1  (j~0  ]rQ1  (h	he]rR1  (hh�eeee]rS1  (hheee]rT1  (j�,  ]rU1  (j�,  ]rV1  (j�,  ]rW1  (h	j�  e]rX1  (hh�e]rY1  (hhe]rZ1  (j�,  ]r[1  (h	h�e]r\1  (hh�e]r]1  (hhe]r^1  (j~0  ]r_1  (h	he]r`1  (hh�eeee]ra1  (hheee]rb1  (j�,  ]rc1  (j�,  ]rd1  (j�,  ]re1  (h	j�  e]rf1  (hh�e]rg1  (hhe]rh1  (j�,  ]ri1  (h	h�e]rj1  (hh�e]rk1  (hhe]rl1  (j~0  ]rm1  (h	he]rn1  (hh�eeee]ro1  (hheeejb1  ]rp1  (j�,  ]rq1  (j�,  ]rr1  (j�,  ]rs1  (h	j�  e]rt1  (hh�e]ru1  (hhe]rv1  (j�,  ]rw1  (h	h�e]rx1  (hh�e]ry1  (hhe]rz1  (j~0  ]r{1  (h	he]r|1  (hh�eeee]r}1  (hheeejp1  jp1  jp1  ]r~1  (j�,  ]r1  (j�,  ]r�1  (j�,  ]r�1  (h	j�  e]r�1  (hh�e]r�1  (hhe]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j~0  ]r�1  (h	he]r�1  (hh�eeee]r�1  (hheeej~1  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (h	j�  e]r�1  (hh�e]r�1  (hhe]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j~0  ]r�1  (h	he]r�1  (hh�eeee]r�1  (hheeej�1  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (h	j�  e]r�1  (hh�e]r�1  (hhe]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j~0  ]r�1  (h	he]r�1  (hh�eeee]r�1  (hheee]r�1  (j�,  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j~0  ]r�1  (h	he]r�1  (hh�eeee]r�1  (hheeej�1  j�1  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j~0  ]r�1  (h	he]r�1  (hh�eeee]r�1  (hheeej�1  j�1  j�1  j�1  j�1  j�1  j�1  j�1  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j~0  ]r�1  (h	he]r�1  (hh�eeee]r�1  (hheee]r�1  (j�,  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j~0  ]r�1  (h	he]r�1  (hh�eeee]r�1  (hheee]r�1  (j�,  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j~0  ]r�1  (h	he]r�1  (hh�eeee]r�1  (hheeej�1  j�1  j�1  j�1  j�1  j�1  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j�,  ]r�1  (h	h�e]r�1  (hh�e]r�1  (hhe]r�1  (j~0  ]r�1  (h	he]r�1  (hh�eeee]r�1  (hheeej�1  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (j�,  ]r�1  (h	h�e]r 2  (hh�e]r2  (hhe]r2  (j�,  ]r2  (h	h�e]r2  (hh�e]r2  (hhe]r2  (j~0  ]r2  (h	he]r2  (hh�eeee]r	2  (hheeej�1  j�1  j�1  j�1  j�1  j�1  j�1  j�1  ]r
2  (j�,  ]r2  (j�,  ]r2  (j�,  ]r2  (h	j�  e]r2  (hh�e]r2  (hhe]r2  (j�,  ]r2  (h	h�e]r2  (hh�e]r2  (hhe]r2  (j~0  ]r2  (h	he]r2  (hh�eeee]r2  (hheee]r2  (j�,  ]r2  (j�,  ]r2  (j�,  ]r2  (h	j�  e]r2  (hh�e]r2  (hhe]r2  (j�,  ]r2  (h	h�e]r 2  (hh�e]r!2  (hhe]r"2  (j~0  ]r#2  (h	he]r$2  (hh�eeee]r%2  (hheeej2  j2  j2  j2  j2  ]r&2  (j�,  ]r'2  (j�,  ]r(2  (j�,  ]r)2  (h	h�e]r*2  (hh�e]r+2  (hhe]r,2  (j�,  ]r-2  (h	h�e]r.2  (hh�e]r/2  (hhe]r02  (j~0  ]r12  (h	he]r22  (hh�eeee]r32  (hheeej&2  j&2  ]r42  (j�,  ]r52  (j�,  ]r62  (j�,  ]r72  (h	h�e]r82  (hh�e]r92  (hhe]r:2  (j�,  ]r;2  (h	h�e]r<2  (hh�e]r=2  (hhe]r>2  (j~0  ]r?2  (h	he]r@2  (hh�eeee]rA2  (hheeej42  j42  j42  j42  j42  j42  j42  ]rB2  (j�,  ]rC2  (j�,  ]rD2  (j�,  ]rE2  (h	h�e]rF2  (hh�e]rG2  (hhe]rH2  (j�,  ]rI2  (h	h�e]rJ2  (hh�e]rK2  (hhe]rL2  (j~0  ]rM2  (h	he]rN2  (hh�eeee]rO2  (hheeejB2  jB2  jB2  jB2  jB2  ]rP2  (j�,  ]rQ2  (j�,  ]rR2  (j�,  ]rS2  (h	h�e]rT2  (hh�e]rU2  (hhe]rV2  (j�,  ]rW2  (h	h�e]rX2  (hh�e]rY2  (hhe]rZ2  (j~0  ]r[2  (h	he]r\2  (hh�eeee]r]2  (hheeejP2  ]r^2  (j�,  ]r_2  (j�,  ]r`2  (j�,  ]ra2  (h	h�e]rb2  (hh�e]rc2  (hhe]rd2  (j�,  ]re2  (h	h�e]rf2  (hh�e]rg2  (hhe]rh2  (j~0  ]ri2  (h	he]rj2  (hh�eeee]rk2  (hheeej^2  ]rl2  (j�,  ]rm2  (j�,  ]rn2  (j�,  ]ro2  (h	h�e]rp2  (hh�e]rq2  (hhe]rr2  (j�,  ]rs2  (h	h�e]rt2  (hh�e]ru2  (hhe]rv2  (j~0  ]rw2  (h	he]rx2  (hh�eeee]ry2  (hheee]rz2  (j�,  ]r{2  (j�,  ]r|2  (j�,  ]r}2  (h	j�  e]r~2  (hh�e]r2  (hhe]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j~0  ]r�2  (h	he]r�2  (hh�eeee]r�2  (hheee]r�2  (j�,  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (h	j�  e]r�2  (hh�e]r�2  (hhe]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j~0  ]r�2  (h	he]r�2  (hh�eeee]r�2  (hheeej�2  j�2  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (h	j�  e]r�2  (hh�e]r�2  (hhe]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j~0  ]r�2  (h	he]r�2  (hh�eeee]r�2  (hheeej�2  j�2  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (h	j�  e]r�2  (hh�e]r�2  (hhe]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j~0  ]r�2  (h	he]r�2  (hh�eeee]r�2  (hheeej�2  j�2  j�2  j�2  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j~0  ]r�2  (h	he]r�2  (hh�eeee]r�2  (hheee]r�2  (j�,  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j~0  ]r�2  (h	he]r�2  (hh�eeee]r�2  (hheeej�2  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j~0  ]r�2  (h	he]r�2  (hh�eeee]r�2  (hheeej�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j~0  ]r�2  (h	he]r�2  (hh�eeee]r�2  (hheeej�2  j�2  j�2  j�2  j�2  j�2  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j~0  ]r�2  (h	he]r�2  (hh�eeee]r�2  (hheeej�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  j�2  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (j�,  ]r�2  (h	h�e]r�2  (hh�e]r�2  (hhe]r�2  (j�,  ]r�2  (h	h�e]r 3  (hh�e]r3  (hhe]r3  (j~0  ]r3  (h	he]r3  (hh�eeee]r3  (hheee]r3  (j�,  ]r3  (j�,  ]r3  (j�,  ]r	3  (h	j�  e]r
3  (hh�e]r3  (hhe]r3  (j�,  ]r3  (h	h�e]r3  (hh�e]r3  (hhe]r3  (j~0  ]r3  (h	he]r3  (hh�eeee]r3  (hheeej3  j3  j3  j3  ]r3  (j�,  ]r3  (j�,  ]r3  (j�,  ]r3  (h	j�  e]r3  (hh�e]r3  (hhe]r3  (j�,  ]r3  (h	h�e]r3  (hh�e]r3  (hhe]r3  (j~0  ]r3  (h	he]r 3  (hh�eeee]r!3  (hheeej3  j3  ]r"3  (j�,  ]r#3  (j�,  ]r$3  (j�,  ]r%3  (h	j�  e]r&3  (hh�e]r'3  (hhe]r(3  (j�,  ]r)3  (h	h�e]r*3  (hh�e]r+3  (hhe]r,3  (j~0  ]r-3  (h	he]r.3  (hh�eeee]r/3  (hheeej"3  j"3  ]r03  (j�,  ]r13  (j�,  ]r23  (j�,  ]r33  (h	j�  e]r43  (hh�e]r53  (hhe]r63  (j�,  ]r73  (h	h�e]r83  (hh�e]r93  (hhe]r:3  (j~0  ]r;3  (h	he]r<3  (hh�eeee]r=3  (hheeej03  j03  j03  j03  ]r>3  (j�,  ]r?3  (j�,  ]r@3  (j�,  ]rA3  (h	j�  e]rB3  (hh�e]rC3  (hhe]rD3  (j�,  ]rE3  (h	h�e]rF3  (hh�e]rG3  (hhe]rH3  (j~0  ]rI3  (h	h�e]rJ3  (hh�eeee]rK3  (hheeej>3  j>3  j>3  j>3  j>3  j>3  j>3  ]rL3  (j�,  ]rM3  (j�,  ]rN3  (j�,  ]rO3  (h	j�  e]rP3  (hh�e]rQ3  (hhe]rR3  (j�,  ]rS3  (h	h�e]rT3  (hh�e]rU3  (hhe]rV3  (j~0  ]rW3  (h	h�e]rX3  (hh�eeee]rY3  (hheeejL3  jL3  ]rZ3  (j�,  ]r[3  (j�,  ]r\3  (j�,  ]r]3  (h	j�  e]r^3  (hh�e]r_3  (hhe]r`3  (j�,  ]ra3  (h	h�e]rb3  (hh�e]rc3  (hhe]rd3  (j~0  ]re3  (h	h�e]rf3  (hh�eeee]rg3  (hheeejZ3  ]rh3  (j�,  ]ri3  (j�,  ]rj3  (j�,  ]rk3  (h	j�  e]rl3  (hh�e]rm3  (hhe]rn3  (j�,  ]ro3  (h	h�e]rp3  (hh�e]rq3  (hhe]rr3  (j~0  ]rs3  (h	h�e]rt3  (hh�eeee]ru3  (hheeejh3  ]rv3  (j�,  ]rw3  (j�,  ]rx3  (j�,  ]ry3  (h	j�  e]rz3  (hh�e]r{3  (hhe]r|3  (j�,  ]r}3  (h	h�e]r~3  (hh�e]r3  (hhe]r�3  (j~0  ]r�3  (h	he]r�3  (hh�eeee]r�3  (hheeejv3  jv3  jv3  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (h	j�  e]r�3  (hh�e]r�3  (hhe]r�3  (j�,  ]r�3  (h	h�e]r�3  (hh�e]r�3  (hhe]r�3  (j~0  ]r�3  (h	he]r�3  (hh�eeee]r�3  (hheeej�3  j�3  j�3  j�3  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (h	j�  e]r�3  (hh�e]r�3  (hhe]r�3  (j�,  ]r�3  (h	h�e]r�3  (hh�e]r�3  (hhe]r�3  (j~0  ]r�3  (h	he]r�3  (hh�eeee]r�3  (hheeej�3  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (h	j�  e]r�3  (hh�e]r�3  (hhe]r�3  (j�,  ]r�3  (h	h�e]r�3  (hh�e]r�3  (hhe]r�3  (j~0  ]r�3  (h	h�e]r�3  (hh�eeee]r�3  (hheeej�3  j�3  j�3  j�3  j�3  j�3  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (h	j�  e]r�3  (hh�e]r�3  (hhe]r�3  (j�,  ]r�3  (h	h�e]r�3  (hh�e]r�3  (hhe]r�3  (j~0  ]r�3  (h	h�e]r�3  (hh�eeee]r�3  (hheeej�3  j�3  j�3  j�3  j�3  j�3  j�3  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (h	j�  e]r�3  (hh�e]r�3  (hhe]r�3  (j�,  ]r�3  (h	h�e]r�3  (hh�e]r�3  (hhe]r�3  (j~0  ]r�3  (h	h�e]r�3  (hh�eeee]r�3  (hheeej�3  j�3  j�3  j�3  j�3  j�3  j�3  j�3  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (h	j�  e]r�3  (hh�e]r�3  (hhe]r�3  (j�,  ]r�3  (h	h�e]r�3  (hh�e]r�3  (hhe]r�3  (j~0  ]r�3  (h	h�e]r�3  (hh�eeee]r�3  (hheeej�3  j�3  j�3  j�3  j�3  j�3  j�3  j�3  j�3  j�3  j�3  j�3  j�3  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (h	j�  e]r�3  (hh�e]r�3  (hhe]r�3  (j�,  ]r�3  (h	h�e]r�3  (hh�e]r�3  (hhe]r�3  (j~0  ]r�3  (h	h�e]r�3  (hh�eeee]r�3  (hheeej�3  j�3  j�3  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (h	j�  e]r�3  (hh�e]r�3  (hhe]r�3  (j�,  ]r�3  (h	h�e]r�3  (hh�e]r�3  (hhe]r�3  (j~0  ]r�3  (h	h�e]r�3  (hh�eeee]r�3  (hheeej�3  j�3  j�3  j�3  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (j�,  ]r�3  (h	j�  e]r�3  (hh�e]r�3  (hhe]r�3  (j�,  ]r�3  (h	h�e]r�3  (hh�e]r�3  (hhe]r�3  (j~0  ]r�3  (h	h�e]r 4  (hh�eeee]r4  (hheee]r4  (j�,  ]r4  (j�,  ]r4  (j�,  ]r4  (h	j�  e]r4  (hh�e]r4  (hhe]r4  (j�,  ]r	4  (h	h�e]r
4  (hh�e]r4  (hhe]r4  (j~0  ]r4  (h	h�e]r4  (hh�eeee]r4  (hheeej4  j4  j4  j4  j4  ]r4  (j�,  ]r4  (j�,  ]r4  (j�,  ]r4  (h	j�  e]r4  (hh�e]r4  (hhe]r4  (j�,  ]r4  (h	h�e]r4  (hh�e]r4  (hhe]r4  (j~0  ]r4  (h	h�e]r4  (hh�eeee]r4  (hheeej4  j4  j4  j4  j4  j4  j4  j4  j4  j4  j4  ]r4  (j�,  ]r4  (j�,  ]r 4  (j�,  ]r!4  (h	j�  e]r"4  (hh�e]r#4  (hhe]r$4  (j�,  ]r%4  (h	h�e]r&4  (hh�e]r'4  (hhe]r(4  (j~0  ]r)4  (h	h�e]r*4  (hh�eeee]r+4  (hheeej4  j4  ]r,4  (j�,  ]r-4  (j�,  ]r.4  (j�,  ]r/4  (h	j�  e]r04  (hh�e]r14  (hhe]r24  (j�,  ]r34  (h	h�e]r44  (hh�e]r54  (hhe]r64  (j~0  ]r74  (h	he]r84  (hh�eeee]r94  (hheeej,4  j,4  j,4  j,4  j,4  ]r:4  (j�,  ]r;4  (j�,  ]r<4  (j�,  ]r=4  (h	j�  e]r>4  (hh�e]r?4  (hhe]r@4  (j�,  ]rA4  (h	h�e]rB4  (hh�e]rC4  (hhe]rD4  (j~0  ]rE4  (h	he]rF4  (hh�eeee]rG4  (hheeej:4  ]rH4  (j�,  ]rI4  (j�,  ]rJ4  (j�,  ]rK4  (h	j�  e]rL4  (hh�e]rM4  (hhe]rN4  (j�,  ]rO4  (h	h�e]rP4  (hh�e]rQ4  (hhe]rR4  (j~0  ]rS4  (h	he]rT4  (hh�eeee]rU4  (hheeejH4  ]rV4  (j�,  ]rW4  (j�,  ]rX4  (j�,  ]rY4  (h	j�  e]rZ4  (hh�e]r[4  (hhe]r\4  (j�,  ]r]4  (h	h�e]r^4  (hh�e]r_4  (hhe]r`4  (j~0  ]ra4  (h	h�e]rb4  (hh�eeee]rc4  (hheeejV4  jV4  jV4  jV4  ]rd4  (j�,  ]re4  (j�,  ]rf4  (j�,  ]rg4  (h	j�  e]rh4  (hh�e]ri4  (hhe]rj4  (j�,  ]rk4  (h	h�e]rl4  (hh�e]rm4  (hhe]rn4  (j~0  ]ro4  (h	he]rp4  (hh�eeee]rq4  (hheeejd4  jd4  jd4  jd4  jd4  jd4  jd4  ]rr4  (j�,  ]rs4  (j�,  ]rt4  (j�,  ]ru4  (h	j�  e]rv4  (hh�e]rw4  (hhe]rx4  (j�,  ]ry4  (h	h�e]rz4  (hh�e]r{4  (hhe]r|4  (j~0  ]r}4  (h	he]r~4  (hh�eeee]r4  (hheeejr4  jr4  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (h	j�  e]r�4  (hh�e]r�4  (hhe]r�4  (j�,  ]r�4  (h	h�e]r�4  (hh�e]r�4  (hhe]r�4  (j~0  ]r�4  (h	he]r�4  (hh�eeee]r�4  (hheeej�4  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (h	j�  e]r�4  (hh�e]r�4  (hhe]r�4  (j�,  ]r�4  (h	h�e]r�4  (hh�e]r�4  (hhe]r�4  (j~0  ]r�4  (h	he]r�4  (hh�eeee]r�4  (hheee]r�4  (j�,  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (h	j�  e]r�4  (hh�e]r�4  (hhe]r�4  (j�,  ]r�4  (h	h�e]r�4  (hh�e]r�4  (hhe]r�4  (j~0  ]r�4  (h	he]r�4  (hh�eeee]r�4  (hheeej�4  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (h	j�  e]r�4  (hh�e]r�4  (hhe]r�4  (j�,  ]r�4  (h	h�e]r�4  (hh�e]r�4  (hhe]r�4  (j~0  ]r�4  (h	he]r�4  (hh�eeee]r�4  (hheee]r�4  (j�,  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (h	j�  e]r�4  (hh�e]r�4  (hhe]r�4  (j�,  ]r�4  (h	h�e]r�4  (hh�e]r�4  (hhe]r�4  (j~0  ]r�4  (h	he]r�4  (hh�eeee]r�4  (hheeej�4  j�4  j�4  j�4  j�4  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (h	j�  e]r�4  (hh�e]r�4  (hhe]r�4  (j�,  ]r�4  (h	h�e]r�4  (hh�e]r�4  (hhe]r�4  (j~0  ]r�4  (h	he]r�4  (hh�eeee]r�4  (hheeej�4  j�4  j�4  j�4  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (h	j�  e]r�4  (hh�e]r�4  (hhe]r�4  (j�,  ]r�4  (h	h�e]r�4  (hh�e]r�4  (hhe]r�4  (j~0  ]r�4  (h	he]r�4  (hh�eeee]r�4  (hheee]r�4  (j�,  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (h	j�  e]r�4  (hh�e]r�4  (hhe]r�4  (j�,  ]r�4  (h	h�e]r�4  (hh�e]r�4  (hhe]r�4  (j~0  ]r�4  (h	h�e]r�4  (hh�eeee]r�4  (hheee]r�4  (j�,  ]r�4  (j�,  ]r�4  (j�,  ]r�4  (h	j�  e]r�4  (hh�e]r�4  (hhe]r�4  (j�,  ]r�4  (h	h�e]r�4  (hh�e]r�4  (hhe]r�4  (j~0  ]r�4  (h	h�e]r�4  (hh�eeee]r�4  (hheeej�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  j�4  ]r�4  (j�,  ]r�4  (j�,  ]r 5  (j�,  ]r5  (h	j�  e]r5  (hh�e]r5  (hhe]r5  (j�,  ]r5  (h	h�e]r5  (hh�e]r5  (hhe]r5  (j~0  ]r	5  (h	h�e]r
5  (hh�eeee]r5  (hheeej�4  j�4  j�4  ]r5  (j�,  ]r5  (j�,  ]r5  (j�,  ]r5  (h	j�  e]r5  (hh�e]r5  (hhe]r5  (j�,  ]r5  (h	h�e]r5  (hh�e]r5  (hhe]r5  (j~0  ]r5  (h	h�e]r5  (hh�eeee]r5  (hheeej5  j5  j5  ]r5  (j�,  ]r5  (j�,  ]r5  (j�,  ]r5  (h	j�  e]r5  (hh�e]r5  (hhe]r 5  (j�,  ]r!5  (h	h�e]r"5  (hh�e]r#5  (hhe]r$5  (j~0  ]r%5  (h	h�e]r&5  (hh�eeee]r'5  (hheee]r(5  (j�,  ]r)5  (j�,  ]r*5  (j�,  ]r+5  (h	j�  e]r,5  (hh�e]r-5  (hhe]r.5  (j�,  ]r/5  (h	h�e]r05  (hh�e]r15  (hhe]r25  (j~0  ]r35  (h	h�e]r45  (hh�eeee]r55  (hheeej(5  j(5  j(5  j(5  j(5  ]r65  (j�,  ]r75  (j�,  ]r85  (j�,  ]r95  (h	j�  e]r:5  (hh�e]r;5  (hhe]r<5  (j�,  ]r=5  (h	h�e]r>5  (hh�e]r?5  (hhe]r@5  (j~0  ]rA5  (h	h�e]rB5  (hh�eeee]rC5  (hheeej65  j65  j65  j65  ]rD5  (j�,  ]rE5  (j�,  ]rF5  (j�,  ]rG5  (h	j�  e]rH5  (hh�e]rI5  (hhe]rJ5  (j�,  ]rK5  (h	h�e]rL5  (hh�e]rM5  (hhe]rN5  (j~0  ]rO5  (h	h�e]rP5  (hh�eeee]rQ5  (hheeejD5  jD5  jD5  jD5  ]rR5  (j�,  ]rS5  (j�,  ]rT5  (j�,  ]rU5  (h	j�  e]rV5  (hh�e]rW5  (hhe]rX5  (j�,  ]rY5  (h	h�e]rZ5  (hh�e]r[5  (hhe]r\5  (j~0  ]r]5  (h	h�e]r^5  (hh�eeee]r_5  (hheee]r`5  (j�,  ]ra5  (j�,  ]rb5  (j�,  ]rc5  (h	j�  e]rd5  (hh�e]re5  (hhe]rf5  (j�,  ]rg5  (h	h�e]rh5  (hh�e]ri5  (hhe]rj5  (j~0  ]rk5  (h	h�e]rl5  (hh�eeee]rm5  (hheee]rn5  (j�,  ]ro5  (j�,  ]rp5  (j�,  ]rq5  (h	j�  e]rr5  (hh�e]rs5  (hhe]rt5  (j�,  ]ru5  (h	h�e]rv5  (hh�e]rw5  (hhe]rx5  (j~0  ]ry5  (h	h�e]rz5  (hh�eeee]r{5  (hheeejn5  jn5  jn5  ]r|5  (j�,  ]r}5  (j�,  ]r~5  (j�,  ]r5  (h	j�  e]r�5  (hh�e]r�5  (hhe]r�5  (j�,  ]r�5  (h	h�e]r�5  (hh�e]r�5  (hhe]r�5  (j~0  ]r�5  (h	h�e]r�5  (hh�eeee]r�5  (hheeej|5  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (h	j�  e]r�5  (hh�e]r�5  (hhe]r�5  (j�,  ]r�5  (h	h�e]r�5  (hh�e]r�5  (hhe]r�5  (j~0  ]r�5  (h	h�e]r�5  (hh�eeee]r�5  (hheee]r�5  (j�,  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (h	j�  e]r�5  (hh�e]r�5  (hhe]r�5  (j�,  ]r�5  (h	h�e]r�5  (hh�e]r�5  (hhe]r�5  (j~0  ]r�5  (h	h�e]r�5  (hh�eeee]r�5  (hheeej�5  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (h	j�  e]r�5  (hh�e]r�5  (hhe]r�5  (j�,  ]r�5  (h	h�e]r�5  (hh�e]r�5  (hhe]r�5  (j~0  ]r�5  (h	h�e]r�5  (hh�eeee]r�5  (hheeej�5  j�5  j�5  j�5  j�5  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (h	j�  e]r�5  (hh�e]r�5  (hhe]r�5  (j�,  ]r�5  (h	h�e]r�5  (hh�e]r�5  (hhe]r�5  (j~0  ]r�5  (h	h�e]r�5  (hh�eeee]r�5  (hheeej�5  j�5  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (h	j�  e]r�5  (hh�e]r�5  (hhe]r�5  (j�,  ]r�5  (h	h�e]r�5  (hh�e]r�5  (hhe]r�5  (j~0  ]r�5  (h	h�e]r�5  (hh�eeee]r�5  (hheee]r�5  (j�,  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (h	j�  e]r�5  (hh�e]r�5  (hhe]r�5  (j�,  ]r�5  (h	h�e]r�5  (hh�e]r�5  (hhe]r�5  (j~0  ]r�5  (h	h�e]r�5  (hh�eeee]r�5  (hheee]r�5  (j�,  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (h	j�  e]r�5  (hh�e]r�5  (hhe]r�5  (j�,  ]r�5  (h	h�e]r�5  (hh�e]r�5  (hhe]r�5  (j~0  ]r�5  (h	h�e]r�5  (hh�eeee]r�5  (hheeej�5  j�5  j�5  j�5  j�5  j�5  j�5  j�5  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (h	j�  e]r�5  (hh�e]r�5  (hhe]r�5  (j�,  ]r�5  (h	h�e]r�5  (hh�e]r�5  (hhe]r�5  (j~0  ]r�5  (h	h�e]r�5  (hh�eeee]r�5  (hheeej�5  j�5  j�5  j�5  j�5  j�5  j�5  j�5  j�5  j�5  j�5  j�5  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (j�,  ]r�5  (h	j�  e]r�5  (hh�e]r�5  (hhe]r 6  (j�,  ]r6  (h	h�e]r6  (hh�e]r6  (hhe]r6  (j~0  ]r6  (h	h�e]r6  (hh�eeee]r6  (hheeej�5  j�5  j�5  j�5  j�5  j�5  j�5  j�5  j�5  ]r6  (j�,  ]r	6  (j�,  ]r
6  (j�,  ]r6  (h	j�  e]r6  (hh�e]r6  (hhe]r6  (j�,  ]r6  (h	h�e]r6  (hh�e]r6  (hhe]r6  (j~0  ]r6  (h	h�e]r6  (hh�eeee]r6  (hheeej6  ]r6  (j�,  ]r6  (j�,  ]r6  (j�,  ]r6  (h	j�  e]r6  (hh�e]r6  (hhe]r6  (j�,  ]r6  (h	h�e]r6  (hh�e]r6  (hhe]r 6  (j~0  ]r!6  (h	h�e]r"6  (hh�eeee]r#6  (hheeej6  j6  j6  j6  ]r$6  (j�,  ]r%6  (j�,  ]r&6  (j�,  ]r'6  (h	j�  e]r(6  (hh�e]r)6  (hhe]r*6  (j�,  ]r+6  (h	h�e]r,6  (hh�e]r-6  (hhe]r.6  (j~0  ]r/6  (h	h�e]r06  (hh�eeee]r16  (hheeej$6  ]r26  (j�,  ]r36  (j�,  ]r46  (j�,  ]r56  (h	j�  e]r66  (hh�e]r76  (hhe]r86  (j�,  ]r96  (h	h�e]r:6  (hh�e]r;6  (hhe]r<6  (j~0  ]r=6  (h	h�e]r>6  (hh�eeee]r?6  (hheeej26  ]r@6  (j�,  ]rA6  (j�,  ]rB6  (j�,  ]rC6  (h	j�  e]rD6  (hh�e]rE6  (hhe]rF6  (j�,  ]rG6  (h	h�e]rH6  (hh�e]rI6  (hhe]rJ6  (j~0  ]rK6  (h	he]rL6  (hh�eeee]rM6  (hheeej@6  j@6  ]rN6  (j�,  ]rO6  (j�,  ]rP6  (j�,  ]rQ6  (h	j�  e]rR6  (hh�e]rS6  (hhe]rT6  (j�,  ]rU6  (h	h�e]rV6  (hh�e]rW6  (hhe]rX6  (j~0  ]rY6  (h	he]rZ6  (hh�eeee]r[6  (hheee]r\6  (j�,  ]r]6  (j�,  ]r^6  (j�,  ]r_6  (h	j�  e]r`6  (hh�e]ra6  (hhe]rb6  (j�,  ]rc6  (h	h�e]rd6  (hh�e]re6  (hhe]rf6  (j~0  ]rg6  (h	he]rh6  (hh�eeee]ri6  (hheeej\6  j\6  j\6  j\6  j\6  ]rj6  (j�,  ]rk6  (j�,  ]rl6  (j�,  ]rm6  (h	j�  e]rn6  (hh�e]ro6  (hhe]rp6  (j�,  ]rq6  (h	h�e]rr6  (hh�e]rs6  (hhe]rt6  (j~0  ]ru6  (h	h�e]rv6  (hh�eeee]rw6  (hheee]rx6  (j�,  ]ry6  (j�,  ]rz6  (j�,  ]r{6  (h	j�  e]r|6  (hh�e]r}6  (hhe]r~6  (j�,  ]r6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j~0  ]r�6  (h	h�e]r�6  (hh�eeee]r�6  (hheeejx6  jx6  jx6  jx6  jx6  jx6  jx6  jx6  jx6  jx6  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (h	j�  e]r�6  (hh�e]r�6  (hhe]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j~0  ]r�6  (h	he]r�6  (hh�eeee]r�6  (hheee]r�6  (j�,  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (h	j�  e]r�6  (hh�e]r�6  (hhe]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j~0  ]r�6  (h	he]r�6  (hh�eeee]r�6  (hheeej�6  j�6  j�6  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j~0  ]r�6  (h	he]r�6  (hh�eeee]r�6  (hheeej�6  j�6  j�6  j�6  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j~0  ]r�6  (h	he]r�6  (hh�eeee]r�6  (hheee]r�6  (j�,  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j~0  ]r�6  (h	he]r�6  (hh�eeee]r�6  (hheee]r�6  (j�,  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j~0  ]r�6  (h	he]r�6  (hh�eeee]r�6  (hheee]r�6  (j�,  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j~0  ]r�6  (h	he]r�6  (hh�eeee]r�6  (hheeej�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j~0  ]r�6  (h	he]r�6  (hh�eeee]r�6  (hheee]r�6  (j�,  ]r�6  (j�,  ]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r�6  (j�,  ]r�6  (h	h�e]r�6  (hh�e]r�6  (hhe]r 7  (j~0  ]r7  (h	he]r7  (hh�eeee]r7  (hheeej�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  j�6  ]r7  (j�,  ]r7  (j�,  ]r7  (j�,  ]r7  (h	h�e]r7  (hh�e]r	7  (hhe]r
7  (j�,  ]r7  (h	h�e]r7  (hh�e]r7  (hhe]r7  (j~0  ]r7  (h	he]r7  (hh�eeee]r7  (hheeej7  j7  ]r7  (j�,  ]r7  (j�,  ]r7  (j�,  ]r7  (h	h�e]r7  (hh�e]r7  (hhe]r7  (j�,  ]r7  (h	h�e]r7  (hh�e]r7  (hhe]r7  (j~0  ]r7  (h	he]r7  (hh�eeee]r7  (hheeej7  j7  ]r 7  (j�,  ]r!7  (j�,  ]r"7  (j�,  ]r#7  (h	h�e]r$7  (hh�e]r%7  (hhe]r&7  (j�,  ]r'7  (h	h�e]r(7  (hh�e]r)7  (hhe]r*7  (j~0  ]r+7  (h	he]r,7  (hh�eeee]r-7  (hheee]r.7  (j�,  ]r/7  (j�,  ]r07  (j�,  ]r17  (h	h�e]r27  (hh�e]r37  (hhe]r47  (j�,  ]r57  (h	h�e]r67  (hh�e]r77  (hhe]r87  (X	   Next-Mover97  ]r:7  (h	he]r;7  (hh�eeee]r<7  (hheeej.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  j.7  ]r=7  (j�,  ]r>7  (j�,  ]r?7  (j�,  ]r@7  (h	h�e]rA7  (hh�e]rB7  (hhe]rC7  (j�,  ]rD7  (h	h�e]rE7  (hh�e]rF7  (hhe]rG7  (j97  ]rH7  (h	he]rI7  (hh�eeee]rJ7  (hheee]rK7  (j�,  ]rL7  (j�,  ]rM7  (j�,  ]rN7  (h	h�e]rO7  (hh�e]rP7  (hhe]rQ7  (j�,  ]rR7  (h	h�e]rS7  (hh�e]rT7  (hhe]rU7  (j97  ]rV7  (h	he]rW7  (hh�eeee]rX7  (hheeejK7  ]rY7  (j�,  ]rZ7  (j�,  ]r[7  (j�,  ]r\7  (h	j�  e]r]7  (hh�e]r^7  (hhe]r_7  (j�,  ]r`7  (h	h�e]ra7  (hh�e]rb7  (hhe]rc7  (j97  ]rd7  (h	he]re7  (hh�eeee]rf7  (hheeejY7  jY7  jY7  ]rg7  (j�,  ]rh7  (j�,  ]ri7  (j�,  ]rj7  (h	j�  e]rk7  (hh�e]rl7  (hhe]rm7  (j�,  ]rn7  (h	h�e]ro7  (hh�e]rp7  (hhe]rq7  (j97  ]rr7  (h	h�e]rs7  (hh�eeee]rt7  (hheee]ru7  (j�,  ]rv7  (j�,  ]rw7  (j�,  ]rx7  (h	j�  e]ry7  (hh�e]rz7  (hhe]r{7  (j�,  ]r|7  (h	h�e]r}7  (hh�e]r~7  (hhe]r7  (j97  ]r�7  (h	h�e]r�7  (hh�eeee]r�7  (hheeeju7  ju7  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (h	j�  e]r�7  (hh�e]r�7  (hhe]r�7  (j�,  ]r�7  (h	h�e]r�7  (hh�e]r�7  (hhe]r�7  (j97  ]r�7  (h	h�e]r�7  (hh�eeee]r�7  (hheee]r�7  (j�,  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (h	j�  e]r�7  (hh�e]r�7  (hhe]r�7  (j�,  ]r�7  (h	h�e]r�7  (hh�e]r�7  (hhe]r�7  (j97  ]r�7  (h	h�e]r�7  (hh�eeee]r�7  (hheeej�7  j�7  j�7  j�7  j�7  j�7  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (h	j�  e]r�7  (hh�e]r�7  (hhe]r�7  (j�,  ]r�7  (h	h�e]r�7  (hh�e]r�7  (hhe]r�7  (j97  ]r�7  (h	h�e]r�7  (hh�eeee]r�7  (hheeej�7  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (h	j�  e]r�7  (hh�e]r�7  (hhe]r�7  (j�,  ]r�7  (h	h�e]r�7  (hh�e]r�7  (hhe]r�7  (j97  ]r�7  (h	h�e]r�7  (hh�eeee]r�7  (hheeej�7  j�7  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (h	j�  e]r�7  (hh�e]r�7  (hhe]r�7  (j�,  ]r�7  (h	h�e]r�7  (hh�e]r�7  (hhe]r�7  (j97  ]r�7  (h	h�e]r�7  (hh�eeee]r�7  (hheeej�7  j�7  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (h	j�  e]r�7  (hh�e]r�7  (hhe]r�7  (j�,  ]r�7  (h	h�e]r�7  (hh�e]r�7  (hhe]r�7  (j97  ]r�7  (h	h�e]r�7  (hh�eeee]r�7  (hheeej�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  j�7  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (h	j�  e]r�7  (hh�e]r�7  (hhe]r�7  (j�,  ]r�7  (h	h�e]r�7  (hh�e]r�7  (hhe]r�7  (j97  ]r�7  (h	he]r�7  (hh�eeee]r�7  (hheeej�7  j�7  j�7  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (h	j�  e]r�7  (hh�e]r�7  (hhe]r�7  (j�,  ]r�7  (h	h�e]r�7  (hh�e]r�7  (hhe]r�7  (j97  ]r�7  (h	he]r�7  (hh�eeee]r�7  (hheee]r�7  (j�,  ]r�7  (j�,  ]r�7  (j�,  ]r�7  (h	j�  e]r�7  (hh�e]r�7  (hhe]r�7  (j�,  ]r�7  (h	h�e]r�7  (hh�e]r�7  (hhe]r�7  (j97  ]r�7  (h	he]r�7  (hh�eeee]r 8  (hheeej�7  ]r8  (j�,  ]r8  (j�,  ]r8  (j�,  ]r8  (h	h�e]r8  (hh�e]r8  (hhe]r8  (j�,  ]r8  (h	h�e]r	8  (hh�e]r
8  (hhe]r8  (j97  ]r8  (h	he]r8  (hh�eeee]r8  (hheee]r8  (j�,  ]r8  (j�,  ]r8  (j�,  ]r8  (h	h�e]r8  (hh�e]r8  (hhe]r8  (j�,  ]r8  (h	h�e]r8  (hh�e]r8  (hhe]r8  (j97  ]r8  (h	he]r8  (hh�eeee]r8  (hheeej8  j8  j8  j8  j8  j8  ]r8  (j�,  ]r8  (j�,  ]r8  (j�,  ]r 8  (h	h�e]r!8  (hh�e]r"8  (hhe]r#8  (j�,  ]r$8  (h	h�e]r%8  (hh�e]r&8  (hhe]r'8  (j97  ]r(8  (h	he]r)8  (hh�eeee]r*8  (hheeej8  ]r+8  (j�,  ]r,8  (j�,  ]r-8  (j�,  ]r.8  (h	h�e]r/8  (hh�e]r08  (hhe]r18  (j�,  ]r28  (h	h�e]r38  (hh�e]r48  (hhe]r58  (j97  ]r68  (h	he]r78  (hh�eeee]r88  (hheeej+8  j+8  j+8  j+8  j+8  j+8  j+8  j+8  j+8  j+8  ]r98  (j�,  ]r:8  (j�,  ]r;8  (j�,  ]r<8  (h	h�e]r=8  (hh�e]r>8  (hhe]r?8  (j�,  ]r@8  (h	h�e]rA8  (hh�e]rB8  (hhe]rC8  (j97  ]rD8  (h	he]rE8  (hh�eeee]rF8  (hheeej98  j98  j98  j98  j98  j98  ]rG8  (j�,  ]rH8  (j�,  ]rI8  (j�,  ]rJ8  (h	h�e]rK8  (hh�e]rL8  (hhe]rM8  (j�,  ]rN8  (h	h�e]rO8  (hh�e]rP8  (hhe]rQ8  (j97  ]rR8  (h	he]rS8  (hh�eeee]rT8  (hheeejG8  jG8  jG8  jG8  jG8  jG8  jG8  jG8  jG8  jG8  jG8  ]rU8  (j�,  ]rV8  (j�,  ]rW8  (j�,  ]rX8  (h	h�e]rY8  (hh�e]rZ8  (hhe]r[8  (j�,  ]r\8  (h	h�e]r]8  (hh�e]r^8  (hhe]r_8  (j97  ]r`8  (h	he]ra8  (hh�eeee]rb8  (hheee]rc8  (j�,  ]rd8  (j�,  ]re8  (j�,  ]rf8  (h	h�e]rg8  (hh�e]rh8  (hhe]ri8  (j�,  ]rj8  (h	h�e]rk8  (hh�e]rl8  (hhe]rm8  (j97  ]rn8  (h	he]ro8  (hh�eeee]rp8  (hheeejc8  jc8  ]rq8  (j�,  ]rr8  (j�,  ]rs8  (j�,  ]rt8  (h	h�e]ru8  (hh�e]rv8  (hhe]rw8  (j�,  ]rx8  (h	h�e]ry8  (hh�e]rz8  (hhe]r{8  (j97  ]r|8  (h	he]r}8  (hh�eeee]r~8  (hheee]r8  (j�,  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j97  ]r�8  (h	he]r�8  (hh�eeee]r�8  (hheee]r�8  (j�,  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j97  ]r�8  (h	he]r�8  (hh�eeee]r�8  (hheee]r�8  (j�,  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j97  ]r�8  (h	he]r�8  (hh�eeee]r�8  (hheee]r�8  (j�,  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j97  ]r�8  (h	he]r�8  (hh�eeee]r�8  (hheeej�8  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j97  ]r�8  (h	he]r�8  (hh�eeee]r�8  (hheeej�8  j�8  j�8  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j97  ]r�8  (h	he]r�8  (hh�eeee]r�8  (hheeej�8  j�8  j�8  j�8  j�8  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (h	j�  e]r�8  (hh�e]r�8  (hhe]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j97  ]r�8  (h	he]r�8  (hh�eeee]r�8  (hheeej�8  j�8  j�8  j�8  j�8  j�8  j�8  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (h	j�  e]r�8  (hh�e]r�8  (hhe]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j97  ]r�8  (h	he]r�8  (hh�eeee]r�8  (hheeej�8  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (j�,  ]r�8  (h	j�  e]r�8  (hh�e]r�8  (hhe]r�8  (j�,  ]r�8  (h	h�e]r�8  (hh�e]r�8  (hhe]r�8  (j97  ]r�8  (h	he]r�8  (hh�eeee]r�8  (hheee]r�8  (j�,  ]r�8  (j�,  ]r�8  (j�,  ]r 9  (h	j�  e]r9  (hh�e]r9  (hhe]r9  (j�,  ]r9  (h	h�e]r9  (hh�e]r9  (hhe]r9  (j97  ]r9  (h	he]r	9  (hh�eeee]r
9  (hheeej�8  j�8  j�8  j�8  ]r9  (j�,  ]r9  (j�,  ]r9  (j�,  ]r9  (h	h�e]r9  (hh�e]r9  (hhe]r9  (j�,  ]r9  (h	h�e]r9  (hh�e]r9  (hhe]r9  (j97  ]r9  (h	he]r9  (hh�eeee]r9  (hheeej9  j9  j9  j9  j9  j9  ]r9  (j�,  ]r9  (j�,  ]r9  (j�,  ]r9  (h	h�e]r9  (hh�e]r9  (hhe]r9  (j�,  ]r 9  (h	h�e]r!9  (hh�e]r"9  (hhe]r#9  (j97  ]r$9  (h	he]r%9  (hh�eeee]r&9  (hheeej9  j9  j9  j9  j9  ]r'9  (j�,  ]r(9  (j�,  ]r)9  (j�,  ]r*9  (h	h�e]r+9  (hh�e]r,9  (hhe]r-9  (j�,  ]r.9  (h	h�e]r/9  (hh�e]r09  (hhe]r19  (j97  ]r29  (h	he]r39  (hh�eeee]r49  (hheeej'9  j'9  j'9  ]r59  (j�,  ]r69  (j�,  ]r79  (j�,  ]r89  (h	h�e]r99  (hh�e]r:9  (hhe]r;9  (j�,  ]r<9  (h	h�e]r=9  (hh�e]r>9  (hhe]r?9  (j97  ]r@9  (h	he]rA9  (hh�eeee]rB9  (hheee]rC9  (j�,  ]rD9  (j�,  ]rE9  (j�,  ]rF9  (h	h�e]rG9  (hh�e]rH9  (hhe]rI9  (j�,  ]rJ9  (h	h�e]rK9  (hh�e]rL9  (hhe]rM9  (j97  ]rN9  (h	he]rO9  (hh�eeee]rP9  (hheeejC9  jC9  jC9  ]rQ9  (j�,  ]rR9  (j�,  ]rS9  (j�,  ]rT9  (h	h�e]rU9  (hh�e]rV9  (hhe]rW9  (j�,  ]rX9  (h	h�e]rY9  (hh�e]rZ9  (hhe]r[9  (j97  ]r\9  (h	he]r]9  (hh�eeee]r^9  (hheeejQ9  jQ9  jQ9  jQ9  ]r_9  (j�,  ]r`9  (j�,  ]ra9  (j�,  ]rb9  (h	h�e]rc9  (hh�e]rd9  (hhe]re9  (j�,  ]rf9  (h	h�e]rg9  (hh�e]rh9  (hhe]ri9  (j97  ]rj9  (h	he]rk9  (hh�eeee]rl9  (hheeej_9  j_9  ]rm9  (j�,  ]rn9  (j�,  ]ro9  (j�,  ]rp9  (h	h�e]rq9  (hh�e]rr9  (hhe]rs9  (j�,  ]rt9  (h	h�e]ru9  (hh�e]rv9  (hhe]rw9  (j97  ]rx9  (h	he]ry9  (hh�eeee]rz9  (hheeejm9  jm9  jm9  jm9  jm9  ]r{9  (j�,  ]r|9  (j�,  ]r}9  (j�,  ]r~9  (h	h�e]r9  (hh�e]r�9  (hhe]r�9  (j�,  ]r�9  (h	h�e]r�9  (hh�e]r�9  (hhe]r�9  (j97  ]r�9  (h	he]r�9  (hh�eeee]r�9  (hheeej{9  j{9  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (h	j�  e]r�9  (hh�e]r�9  (hhe]r�9  (j�,  ]r�9  (h	h�e]r�9  (hh�e]r�9  (hhe]r�9  (j97  ]r�9  (h	he]r�9  (hh�eeee]r�9  (hheeej�9  j�9  j�9  j�9  j�9  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (h	j�  e]r�9  (hh�e]r�9  (hhe]r�9  (j�,  ]r�9  (h	h�e]r�9  (hh�e]r�9  (hhe]r�9  (j97  ]r�9  (h	he]r�9  (hh�eeee]r�9  (hheeej�9  j�9  j�9  j�9  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (h	j�  e]r�9  (hh�e]r�9  (hhe]r�9  (j�,  ]r�9  (h	h�e]r�9  (hh�e]r�9  (hhe]r�9  (j97  ]r�9  (h	he]r�9  (hh�eeee]r�9  (hheeej�9  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (h	j�  e]r�9  (hh�e]r�9  (hhe]r�9  (j�,  ]r�9  (h	h�e]r�9  (hh�e]r�9  (hhe]r�9  (j97  ]r�9  (h	he]r�9  (hh�eeee]r�9  (hheeej�9  j�9  j�9  j�9  j�9  j�9  j�9  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (h	j�  e]r�9  (hh�e]r�9  (hhe]r�9  (j�,  ]r�9  (h	h�e]r�9  (hh�e]r�9  (hhe]r�9  (j97  ]r�9  (h	he]r�9  (hh�eeee]r�9  (hheeej�9  j�9  j�9  j�9  j�9  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (h	j�  e]r�9  (hh�e]r�9  (hhe]r�9  (j�,  ]r�9  (h	h�e]r�9  (hh�e]r�9  (hhe]r�9  (j97  ]r�9  (h	he]r�9  (hh�eeee]r�9  (hheee]r�9  (j�,  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (h	j�  e]r�9  (hh�e]r�9  (hhe]r�9  (j�,  ]r�9  (h	h�e]r�9  (hh�e]r�9  (hhe]r�9  (j97  ]r�9  (h	he]r�9  (hh�eeee]r�9  (hheeej�9  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (h	j�  e]r�9  (hh�e]r�9  (hhe]r�9  (j�,  ]r�9  (h	h�e]r�9  (hh�e]r�9  (hhe]r�9  (j97  ]r�9  (h	he]r�9  (hh�eeee]r�9  (hheeej�9  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (j�,  ]r�9  (h	j�  e]r�9  (hh�e]r�9  (hhe]r�9  (j�,  ]r :  (h	h�e]r:  (hh�e]r:  (hhe]r:  (j97  ]r:  (h	he]r:  (hh�eeee]r:  (hheee]r:  (j�,  ]r:  (j�,  ]r	:  (j�,  ]r
:  (h	j�  e]r:  (hh�e]r:  (hhe]r:  (j�,  ]r:  (h	h�e]r:  (hh�e]r:  (hhe]r:  (j97  ]r:  (h	he]r:  (hh�eeee]r:  (hheeej:  j:  j:  j:  j:  j:  ]r:  (j�,  ]r:  (j�,  ]r:  (j�,  ]r:  (h	j�  e]r:  (hh�e]r:  (hhe]r:  (j�,  ]r:  (h	h�e]r:  (hh�e]r:  (hhe]r:  (j97  ]r :  (h	he]r!:  (hh�eeee]r":  (hheeej:  j:  ]r#:  (j�,  ]r$:  (j�,  ]r%:  (j�,  ]r&:  (h	h�e]r':  (hh�e]r(:  (hhe]r):  (j�,  ]r*:  (h	h�e]r+:  (hh�e]r,:  (hhe]r-:  (j97  ]r.:  (h	he]r/:  (hh�eeee]r0:  (hheeej#:  ]r1:  (j�,  ]r2:  (j�,  ]r3:  (j�,  ]r4:  (h	h�e]r5:  (hh�e]r6:  (hhe]r7:  (j�,  ]r8:  (h	h�e]r9:  (hh�e]r::  (hhe]r;:  (j97  ]r<:  (h	he]r=:  (hh�eeee]r>:  (hheeej1:  e(j1:  j1:  ]r?:  (j�,  ]r@:  (j�,  ]rA:  (j�,  ]rB:  (h	h�e]rC:  (hh�e]rD:  (hhe]rE:  (j�,  ]rF:  (h	h�e]rG:  (hh�e]rH:  (hhe]rI:  (j97  ]rJ:  (h	he]rK:  (hh�eeee]rL:  (hheeej?:  j?:  j?:  j?:  j?:  j?:  j?:  j?:  j?:  j?:  j?:  j?:  j?:  j?:  j?:  ]rM:  (j�,  ]rN:  (j�,  ]rO:  (j�,  ]rP:  (h	h�e]rQ:  (hh�e]rR:  (hhe]rS:  (j�,  ]rT:  (h	h�e]rU:  (hh�e]rV:  (hhe]rW:  (j97  ]rX:  (h	he]rY:  (hh�eeee]rZ:  (hheee]r[:  (j�,  ]r\:  (j�,  ]r]:  (j�,  ]r^:  (h	h�e]r_:  (hh�e]r`:  (hhe]ra:  (j�,  ]rb:  (h	h�e]rc:  (hh�e]rd:  (hhe]re:  (j97  ]rf:  (h	he]rg:  (hh�eeee]rh:  (hheee]ri:  (j�,  ]rj:  (j�,  ]rk:  (j�,  ]rl:  (h	h�e]rm:  (hh�e]rn:  (hhe]ro:  (j�,  ]rp:  (h	h�e]rq:  (hh�e]rr:  (hhe]rs:  (j97  ]rt:  (h	he]ru:  (hh�eeee]rv:  (hheeeji:  ]rw:  (j�,  ]rx:  (j�,  ]ry:  (j�,  ]rz:  (h	j�  e]r{:  (hh�e]r|:  (hhe]r}:  (j�,  ]r~:  (h	h�e]r:  (hh�e]r�:  (hhe]r�:  (j97  ]r�:  (h	he]r�:  (hh�eeee]r�:  (hheeejw:  jw:  jw:  jw:  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (h	j�  e]r�:  (hh�e]r�:  (hhe]r�:  (j�,  ]r�:  (h	h�e]r�:  (hh�e]r�:  (hhe]r�:  (j97  ]r�:  (h	he]r�:  (hh�eeee]r�:  (hheeej�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (h	j�  e]r�:  (hh�e]r�:  (hhe]r�:  (j�,  ]r�:  (h	h�e]r�:  (hh�e]r�:  (hhe]r�:  (j97  ]r�:  (h	he]r�:  (hh�eeee]r�:  (hheeej�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (h	j�  e]r�:  (hh�e]r�:  (hhe]r�:  (j�,  ]r�:  (h	h�e]r�:  (hh�e]r�:  (hhe]r�:  (j97  ]r�:  (h	he]r�:  (hh�eeee]r�:  (hheeej�:  j�:  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (h	j�  e]r�:  (hh�e]r�:  (hhe]r�:  (j�,  ]r�:  (h	h�e]r�:  (hh�e]r�:  (hhe]r�:  (j97  ]r�:  (h	he]r�:  (hh�eeee]r�:  (hheeej�:  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (h	j�  e]r�:  (hh�e]r�:  (hhe]r�:  (j�,  ]r�:  (h	h�e]r�:  (hh�e]r�:  (hhe]r�:  (j97  ]r�:  (h	he]r�:  (hh�eeee]r�:  (hheeej�:  j�:  j�:  j�:  j�:  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (h	j�  e]r�:  (hh�e]r�:  (hhe]r�:  (j�,  ]r�:  (h	h�e]r�:  (hh�e]r�:  (hhe]r�:  (j97  ]r�:  (h	he]r�:  (hh�eeee]r�:  (hheeej�:  j�:  j�:  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (h	j�  e]r�:  (hh�e]r�:  (hhe]r�:  (j�,  ]r�:  (h	h�e]r�:  (hh�e]r�:  (hhe]r�:  (j97  ]r�:  (h	he]r�:  (hh�eeee]r�:  (hheeej�:  j�:  j�:  j�:  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (h	j�  e]r�:  (hh�e]r�:  (hhe]r�:  (j�,  ]r�:  (h	h�e]r�:  (hh�e]r�:  (hhe]r�:  (j97  ]r�:  (h	he]r�:  (hh�eeee]r�:  (hheeej�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  j�:  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (j�,  ]r�:  (h	j�  e]r�:  (hh�e]r�:  (hhe]r�:  (j�,  ]r�:  (h	h�e]r�:  (hh�e]r�:  (hhe]r�:  (j97  ]r ;  (h	he]r;  (hh�eeee]r;  (hheeej�:  ]r;  (j�,  ]r;  (j�,  ]r;  (j�,  ]r;  (h	j�  e]r;  (hh�e]r;  (hhe]r	;  (j�,  ]r
;  (h	h�e]r;  (hh�e]r;  (hhe]r;  (j97  ]r;  (h	he]r;  (hh�eeee]r;  (hheeej;  j;  ]r;  (j�,  ]r;  (j�,  ]r;  (j�,  ]r;  (h	j�  e]r;  (hh�e]r;  (hhe]r;  (j�,  ]r;  (h	h�e]r;  (hh�e]r;  (hhe]r;  (j97  ]r;  (h	he]r;  (hh�eeee]r;  (hheee]r;  (j�,  ]r ;  (j�,  ]r!;  (j�,  ]r";  (h	j�  e]r#;  (hh�e]r$;  (hhe]r%;  (j�,  ]r&;  (h	h�e]r';  (hh�e]r(;  (hhe]r);  (j97  ]r*;  (h	he]r+;  (hh�eeee]r,;  (hheee]r-;  (j�,  ]r.;  (j�,  ]r/;  (j�,  ]r0;  (h	j�  e]r1;  (hh�e]r2;  (hhe]r3;  (j�,  ]r4;  (h	h�e]r5;  (hh�e]r6;  (hhe]r7;  (j97  ]r8;  (h	he]r9;  (hh�eeee]r:;  (hheeej-;  j-;  j-;  j-;  ]r;;  (j�,  ]r<;  (j�,  ]r=;  (j�,  ]r>;  (h	j�  e]r?;  (hh�e]r@;  (hhe]rA;  (j�,  ]rB;  (h	h�e]rC;  (hh�e]rD;  (hhe]rE;  (j97  ]rF;  (h	he]rG;  (hh�eeee]rH;  (hheeej;;  j;;  j;;  ]rI;  (j�,  ]rJ;  (j�,  ]rK;  (j�,  ]rL;  (h	j�  e]rM;  (hh�e]rN;  (hhe]rO;  (j�,  ]rP;  (h	h�e]rQ;  (hh�e]rR;  (hhe]rS;  (j97  ]rT;  (h	he]rU;  (hh�eeee]rV;  (hheeejI;  jI;  jI;  jI;  jI;  jI;  ]rW;  (j�,  ]rX;  (j�,  ]rY;  (j�,  ]rZ;  (h	j�  e]r[;  (hh�e]r\;  (hhe]r];  (j�,  ]r^;  (h	h�e]r_;  (hh�e]r`;  (hhe]ra;  (j97  ]rb;  (h	he]rc;  (hh�eeee]rd;  (hheeejW;  jW;  jW;  ]re;  (j�,  ]rf;  (j�,  ]rg;  (j�,  ]rh;  (h	j�  e]ri;  (hh�e]rj;  (hhe]rk;  (j�,  ]rl;  (h	h�e]rm;  (hh�e]rn;  (hhe]ro;  (j97  ]rp;  (h	he]rq;  (hh�eeee]rr;  (hheeeje;  je;  ]rs;  (j�,  ]rt;  (j�,  ]ru;  (j�,  ]rv;  (h	j�  e]rw;  (hh�e]rx;  (hhe]ry;  (j�,  ]rz;  (h	h�e]r{;  (hh�e]r|;  (hhe]r};  (j97  ]r~;  (h	he]r;  (hh�eeee]r�;  (hheeejs;  js;  js;  js;  js;  js;  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (h	j�  e]r�;  (hh�e]r�;  (hhe]r�;  (j�,  ]r�;  (h	h�e]r�;  (hh�e]r�;  (hhe]r�;  (j97  ]r�;  (h	he]r�;  (hh�eeee]r�;  (hheeej�;  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (h	j�  e]r�;  (hh�e]r�;  (hhe]r�;  (j�,  ]r�;  (h	h�e]r�;  (hh�e]r�;  (hhe]r�;  (j97  ]r�;  (h	he]r�;  (hh�eeee]r�;  (hheeej�;  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (h	j�  e]r�;  (hh�e]r�;  (hhe]r�;  (j�,  ]r�;  (h	h�e]r�;  (hh�e]r�;  (hhe]r�;  (j97  ]r�;  (h	he]r�;  (hh�eeee]r�;  (hheeej�;  j�;  j�;  j�;  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (h	j�  e]r�;  (hh�e]r�;  (hhe]r�;  (j�,  ]r�;  (h	h�e]r�;  (hh�e]r�;  (hhe]r�;  (j97  ]r�;  (h	he]r�;  (hh�eeee]r�;  (hheeej�;  j�;  j�;  j�;  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (h	j�  e]r�;  (hh�e]r�;  (hhe]r�;  (j�,  ]r�;  (h	h�e]r�;  (hh�e]r�;  (hhe]r�;  (j97  ]r�;  (h	he]r�;  (hh�eeee]r�;  (hheeej�;  j�;  j�;  j�;  j�;  j�;  j�;  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (h	j�  e]r�;  (hh�e]r�;  (hhe]r�;  (j�,  ]r�;  (h	h�e]r�;  (hh�e]r�;  (hhe]r�;  (j97  ]r�;  (h	he]r�;  (hh�eeee]r�;  (hheeej�;  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (h	j�  e]r�;  (hh�e]r�;  (hhe]r�;  (j�,  ]r�;  (h	h�e]r�;  (hh�e]r�;  (hhe]r�;  (j97  ]r�;  (h	he]r�;  (hh�eeee]r�;  (hheeej�;  j�;  j�;  j�;  j�;  j�;  j�;  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (h	j�  e]r�;  (hh�e]r�;  (hhe]r�;  (j�,  ]r�;  (h	h�e]r�;  (hh�e]r�;  (hhe]r�;  (j97  ]r�;  (h	he]r�;  (hh�eeee]r�;  (hheeej�;  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (j�,  ]r�;  (h	j�  e]r�;  (hh�e]r�;  (hhe]r�;  (j�,  ]r�;  (h	h�e]r�;  (hh�e]r�;  (hhe]r�;  (j97  ]r�;  (h	he]r�;  (hh�eeee]r�;  (hheee]r�;  (j�,  ]r <  (j�,  ]r<  (j�,  ]r<  (h	j�  e]r<  (hh�e]r<  (hhe]r<  (j�,  ]r<  (h	h�e]r<  (hh�e]r<  (hhe]r	<  (j97  ]r
<  (h	he]r<  (hh�eeee]r<  (hheee]r<  (j�,  ]r<  (j�,  ]r<  (j�,  ]r<  (h	j�  e]r<  (hh�e]r<  (hhe]r<  (j�,  ]r<  (h	h�e]r<  (hh�e]r<  (hhe]r<  (j97  ]r<  (h	he]r<  (hh�eeee]r<  (hheeej<  j<  j<  ]r<  (j�,  ]r<  (j�,  ]r<  (j�,  ]r<  (h	j�  e]r<  (hh�e]r <  (hhe]r!<  (j�,  ]r"<  (h	h�e]r#<  (hh�e]r$<  (hhe]r%<  (j97  ]r&<  (h	he]r'<  (hh�eeee]r(<  (hheeej<  j<  j<  j<  j<  j<  j<  j<  j<  j<  j<  j<  ]r)<  (j�,  ]r*<  (j�,  ]r+<  (j�,  ]r,<  (h	j�  e]r-<  (hh�e]r.<  (hhe]r/<  (j�,  ]r0<  (h	h�e]r1<  (hh�e]r2<  (hhe]r3<  (j97  ]r4<  (h	he]r5<  (hh�eeee]r6<  (hheee]r7<  (j�,  ]r8<  (j�,  ]r9<  (j�,  ]r:<  (h	j�  e]r;<  (hh�e]r<<  (hhe]r=<  (j�,  ]r><  (h	h�e]r?<  (hh�e]r@<  (hhe]rA<  (j97  ]rB<  (h	he]rC<  (hh�eeee]rD<  (hheeej7<  ]rE<  (j�,  ]rF<  (j�,  ]rG<  (j�,  ]rH<  (h	j�  e]rI<  (hh�e]rJ<  (hhe]rK<  (j�,  ]rL<  (h	h�e]rM<  (hh�e]rN<  (hhe]rO<  (j97  ]rP<  (h	he]rQ<  (hh�eeee]rR<  (hheeejE<  jE<  jE<  ]rS<  (j�,  ]rT<  (j�,  ]rU<  (j�,  ]rV<  (h	j�  e]rW<  (hh�e]rX<  (hhe]rY<  (j�,  ]rZ<  (h	h�e]r[<  (hh�e]r\<  (hhe]r]<  (j97  ]r^<  (h	he]r_<  (hh�eeee]r`<  (hheee]ra<  (j�,  ]rb<  (j�,  ]rc<  (j�,  ]rd<  (h	j�  e]re<  (hh�e]rf<  (hhe]rg<  (j�,  ]rh<  (h	h�e]ri<  (hh�e]rj<  (hhe]rk<  (j97  ]rl<  (h	he]rm<  (hh�eeee]rn<  (hheeeja<  ja<  ja<  ja<  ]ro<  (j�,  ]rp<  (j�,  ]rq<  (j�,  ]rr<  (h	j�  e]rs<  (hh�e]rt<  (hhe]ru<  (j�,  ]rv<  (h	h�e]rw<  (hh�e]rx<  (hhe]ry<  (j97  ]rz<  (h	he]r{<  (hh�eeee]r|<  (hheeejo<  jo<  jo<  jo<  jo<  ]r}<  (j�,  ]r~<  (j�,  ]r<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j97  ]r�<  (h	he]r�<  (hh�eeee]r�<  (hheeej}<  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j97  ]r�<  (h	he]r�<  (hh�eeee]r�<  (hheeej�<  j�<  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j97  ]r�<  (h	he]r�<  (hh�eeee]r�<  (hheeej�<  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j97  ]r�<  (h	he]r�<  (hh�eeee]r�<  (hheeej�<  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j97  ]r�<  (h	he]r�<  (hh�eeee]r�<  (hheeej�<  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j97  ]r�<  (h	he]r�<  (hh�eeee]r�<  (hheee]r�<  (j�,  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j97  ]r�<  (h	he]r�<  (hh�eeee]r�<  (hheee]r�<  (j�,  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j97  ]r�<  (h	he]r�<  (hh�eeee]r�<  (hheeej�<  j�<  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (h	j�  e]r�<  (hh�e]r�<  (hhe]r�<  (j�,  ]r�<  (h	h�e]r�<  (hh�e]r�<  (hhe]r�<  (j97  ]r�<  (h	he]r�<  (hh�eeee]r�<  (hheee]r�<  (j�,  ]r�<  (j�,  ]r�<  (j�,  ]r�<  (h	j�  e]r�<  (hh�e]r =  (hhe]r=  (j�,  ]r=  (h	h�e]r=  (hh�e]r=  (hhe]r=  (j97  ]r=  (h	he]r=  (hh�eeee]r=  (hheeej�<  ]r	=  (j�,  ]r
=  (j�,  ]r=  (j�,  ]r=  (h	j�  e]r=  (hh�e]r=  (hhe]r=  (j�,  ]r=  (h	h�e]r=  (hh�e]r=  (hhe]r=  (j97  ]r=  (h	he]r=  (hh�eeee]r=  (hheeej	=  j	=  j	=  j	=  j	=  ]r=  (j�,  ]r=  (j�,  ]r=  (j�,  ]r=  (h	j�  e]r=  (hh�e]r=  (hhe]r=  (j�,  ]r=  (h	h�e]r=  (hh�e]r =  (hhe]r!=  (j97  ]r"=  (h	he]r#=  (hh�eeee]r$=  (hheeej=  ]r%=  (j�,  ]r&=  (j�,  ]r'=  (j�,  ]r(=  (h	j�  e]r)=  (hh�e]r*=  (hhe]r+=  (j�,  ]r,=  (h	h�e]r-=  (hh�e]r.=  (hhe]r/=  (j97  ]r0=  (h	he]r1=  (hh�eeee]r2=  (hheeej%=  j%=  j%=  j%=  ]r3=  (j�,  ]r4=  (j�,  ]r5=  (j�,  ]r6=  (h	j�  e]r7=  (hh�e]r8=  (hhe]r9=  (j�,  ]r:=  (h	h�e]r;=  (hh�e]r<=  (hhe]r==  (j97  ]r>=  (h	he]r?=  (hh�eeee]r@=  (hheeej3=  j3=  j3=  ]rA=  (j�,  ]rB=  (j�,  ]rC=  (j�,  ]rD=  (h	j�  e]rE=  (hh�e]rF=  (hhe]rG=  (j�,  ]rH=  (h	h�e]rI=  (hh�e]rJ=  (hhe]rK=  (j97  ]rL=  (h	he]rM=  (hh�eeee]rN=  (hheeejA=  ]rO=  (j�,  ]rP=  (j�,  ]rQ=  (j�,  ]rR=  (h	j�  e]rS=  (hh�e]rT=  (hhe]rU=  (j�,  ]rV=  (h	h�e]rW=  (hh�e]rX=  (hhe]rY=  (j97  ]rZ=  (h	he]r[=  (hh�eeee]r\=  (hheeejO=  jO=  ]r]=  (j�,  ]r^=  (j�,  ]r_=  (j�,  ]r`=  (h	j�  e]ra=  (hh�e]rb=  (hhe]rc=  (j�,  ]rd=  (h	h�e]re=  (hh�e]rf=  (hhe]rg=  (j97  ]rh=  (h	he]ri=  (hh�eeee]rj=  (hheeej]=  ]rk=  (j�,  ]rl=  (j�,  ]rm=  (j�,  ]rn=  (h	j�  e]ro=  (hh�e]rp=  (hhe]rq=  (j�,  ]rr=  (h	h�e]rs=  (hh�e]rt=  (hhe]ru=  (j97  ]rv=  (h	he]rw=  (hh�eeee]rx=  (hheeejk=  ]ry=  (j�,  ]rz=  (j�,  ]r{=  (j�,  ]r|=  (h	j�  e]r}=  (hh�e]r~=  (hhe]r=  (j�,  ]r�=  (h	h�e]r�=  (hh�e]r�=  (hhe]r�=  (j97  ]r�=  (h	he]r�=  (hh�eeee]r�=  (hheeejy=  jy=  jy=  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (h	j�  e]r�=  (hh�e]r�=  (hhe]r�=  (j�,  ]r�=  (h	h�e]r�=  (hh�e]r�=  (hhe]r�=  (j97  ]r�=  (h	he]r�=  (hh�eeee]r�=  (hheeej�=  j�=  j�=  j�=  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (h	j�  e]r�=  (hh�e]r�=  (hhe]r�=  (j�,  ]r�=  (h	h�e]r�=  (hh�e]r�=  (hhe]r�=  (j97  ]r�=  (h	he]r�=  (hh�eeee]r�=  (hheeej�=  j�=  j�=  j�=  j�=  j�=  j�=  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (h	j�  e]r�=  (hh�e]r�=  (hhe]r�=  (j�,  ]r�=  (h	h�e]r�=  (hh�e]r�=  (hhe]r�=  (j97  ]r�=  (h	he]r�=  (hh�eeee]r�=  (hheeej�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (h	j�  e]r�=  (hh�e]r�=  (hhe]r�=  (j�,  ]r�=  (h	h�e]r�=  (hh�e]r�=  (hhe]r�=  (j97  ]r�=  (h	he]r�=  (hh�eeee]r�=  (hheeej�=  j�=  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (h	j�  e]r�=  (hh�e]r�=  (hhe]r�=  (j�,  ]r�=  (h	h�e]r�=  (hh�e]r�=  (hhe]r�=  (j97  ]r�=  (h	he]r�=  (hh�eeee]r�=  (hheeej�=  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (h	j�  e]r�=  (hh�e]r�=  (hhe]r�=  (j�,  ]r�=  (h	h�e]r�=  (hh�e]r�=  (hhe]r�=  (j97  ]r�=  (h	he]r�=  (hh�eeee]r�=  (hheeej�=  j�=  j�=  j�=  j�=  j�=  j�=  j�=  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (h	j�  e]r�=  (hh�e]r�=  (hhe]r�=  (j�,  ]r�=  (h	h�e]r�=  (hh�e]r�=  (hhe]r�=  (j97  ]r�=  (h	he]r�=  (hh�eeee]r�=  (hheee]r�=  (j�,  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (h	j�  e]r�=  (hh�e]r�=  (hhe]r�=  (j�,  ]r�=  (h	h�e]r�=  (hh�e]r�=  (hhe]r�=  (j97  ]r�=  (h	he]r�=  (hh�eeee]r�=  (hheeej�=  j�=  j�=  j�=  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (j�,  ]r�=  (h	j�  e]r�=  (hh�e]r�=  (hhe]r�=  (j�,  ]r�=  (h	h�e]r�=  (hh�e]r >  (hhe]r>  (j97  ]r>  (h	he]r>  (hh�eeee]r>  (hheeej�=  ]r>  (j�,  ]r>  (j�,  ]r>  (j�,  ]r>  (h	j�  e]r	>  (hh�e]r
>  (hhe]r>  (j�,  ]r>  (h	h�e]r>  (hh�e]r>  (hhe]r>  (j97  ]r>  (h	he]r>  (hh�eeee]r>  (hheeej>  ]r>  (j�,  ]r>  (j�,  ]r>  (j�,  ]r>  (h	j�  e]r>  (hh�e]r>  (hhe]r>  (j�,  ]r>  (h	h�e]r>  (hh�e]r>  (hhe]r>  (j97  ]r>  (h	he]r>  (hh�eeee]r >  (hheeej>  j>  j>  j>  j>  j>  j>  j>  ]r!>  (j�,  ]r">  (j�,  ]r#>  (j�,  ]r$>  (h	j�  e]r%>  (hh�e]r&>  (hhe]r'>  (j�,  ]r(>  (h	h�e]r)>  (hh�e]r*>  (hhe]r+>  (j97  ]r,>  (h	he]r->  (hh�eeee]r.>  (hheeej!>  j!>  j!>  j!>  j!>  j!>  j!>  j!>  ]r/>  (j�,  ]r0>  (j�,  ]r1>  (j�,  ]r2>  (h	j�  e]r3>  (hh�e]r4>  (hhe]r5>  (j�,  ]r6>  (h	h�e]r7>  (hh�e]r8>  (hhe]r9>  (j97  ]r:>  (h	he]r;>  (hh�eeee]r<>  (hheeej/>  j/>  j/>  j/>  ]r=>  (j�,  ]r>>  (j�,  ]r?>  (j�,  ]r@>  (h	j�  e]rA>  (hh�e]rB>  (hhe]rC>  (X   MovedrD>  ]rE>  (h	he]rF>  (hh�e]rG>  (hhe]rH>  (X	   Next-MoverI>  ]rJ>  (h	h�e]rK>  (hh�eeee]rL>  (hheeej=>  j=>  j=>  j=>  j=>  j=>  j=>  j=>  ]rM>  (j�,  ]rN>  (j�,  ]rO>  (j�,  ]rP>  (h	j�  e]rQ>  (hh�e]rR>  (hhe]rS>  (jD>  ]rT>  (h	he]rU>  (hh�e]rV>  (hhe]rW>  (jI>  ]rX>  (h	h�e]rY>  (hh�eeee]rZ>  (hheeejM>  jM>  jM>  jM>  ]r[>  (j�,  ]r\>  (j�,  ]r]>  (j�,  ]r^>  (h	j�  e]r_>  (hh�e]r`>  (hhe]ra>  (jD>  ]rb>  (h	he]rc>  (hh�e]rd>  (hhe]re>  (jI>  ]rf>  (h	h�e]rg>  (hh�eeee]rh>  (hheeej[>  j[>  j[>  ]ri>  (j�,  ]rj>  (j�,  ]rk>  (j�,  ]rl>  (h	j�  e]rm>  (hh�e]rn>  (hhe]ro>  (jD>  ]rp>  (h	he]rq>  (hh�e]rr>  (hhe]rs>  (jI>  ]rt>  (h	h�e]ru>  (hh�eeee]rv>  (hheee]rw>  (j�,  ]rx>  (j�,  ]ry>  (j�,  ]rz>  (h	h�e]r{>  (hh�e]r|>  (hhe]r}>  (jD>  ]r~>  (h	he]r>  (hh�e]r�>  (hhe]r�>  (jI>  ]r�>  (h	h�e]r�>  (hh�eeee]r�>  (hheeejw>  jw>  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (h	h�e]r�>  (hh�e]r�>  (hhe]r�>  (jD>  ]r�>  (h	he]r�>  (hh�e]r�>  (hhe]r�>  (jI>  ]r�>  (h	h�e]r�>  (hh�eeee]r�>  (hheeej�>  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (h	h�e]r�>  (hh�e]r�>  (hhe]r�>  (jD>  ]r�>  (h	he]r�>  (hh�e]r�>  (hhe]r�>  (jI>  ]r�>  (h	h�e]r�>  (hh�eeee]r�>  (hheeej�>  j�>  j�>  j�>  j�>  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (h	h�e]r�>  (hh�e]r�>  (hhe]r�>  (jD>  ]r�>  (h	he]r�>  (hh�e]r�>  (hhe]r�>  (jI>  ]r�>  (h	h�e]r�>  (hh�eeee]r�>  (hheeej�>  j�>  j�>  j�>  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (h	h�e]r�>  (hh�e]r�>  (hhe]r�>  (jD>  ]r�>  (h	he]r�>  (hh�e]r�>  (hhe]r�>  (jI>  ]r�>  (h	h�e]r�>  (hh�eeee]r�>  (hheee]r�>  (j�,  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (h	h�e]r�>  (hh�e]r�>  (hhe]r�>  (jD>  ]r�>  (h	he]r�>  (hh�e]r�>  (hhe]r�>  (jI>  ]r�>  (h	h�e]r�>  (hh�eeee]r�>  (hheeej�>  j�>  j�>  j�>  j�>  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (h	h�e]r�>  (hh�e]r�>  (hhe]r�>  (jD>  ]r�>  (h	he]r�>  (hh�e]r�>  (hhe]r�>  (jI>  ]r�>  (h	h�e]r�>  (hh�eeee]r�>  (hheeej�>  j�>  j�>  j�>  j�>  j�>  j�>  j�>  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (h	h�e]r�>  (hh�e]r�>  (hhe]r�>  (jD>  ]r�>  (h	he]r�>  (hh�e]r�>  (hhe]r�>  (jI>  ]r�>  (h	h�e]r�>  (hh�eeee]r�>  (hheeej�>  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (h	h�e]r�>  (hh�e]r�>  (hhe]r�>  (jD>  ]r�>  (h	he]r�>  (hh�e]r�>  (hhe]r�>  (jI>  ]r�>  (h	h�e]r�>  (hh�eeee]r�>  (hheee]r�>  (j�,  ]r�>  (j�,  ]r�>  (j�,  ]r�>  (h	h�e]r�>  (hh�e]r�>  (hhe]r�>  (jD>  ]r�>  (h	he]r�>  (hh�e]r�>  (hhe]r�>  (jI>  ]r ?  (h	h�e]r?  (hh�eeee]r?  (hheeej�>  j�>  j�>  j�>  j�>  j�>  j�>  j�>  ]r?  (j�,  ]r?  (j�,  ]r?  (j�,  ]r?  (h	h�e]r?  (hh�e]r?  (hhe]r	?  (jD>  ]r
?  (h	he]r?  (hh�e]r?  (hhe]r?  (jI>  ]r?  (h	h�e]r?  (hh�eeee]r?  (hheeej?  j?  j?  j?  j?  ]r?  (j�,  ]r?  (j�,  ]r?  (j�,  ]r?  (h	h�e]r?  (hh�e]r?  (hhe]r?  (jD>  ]r?  (h	he]r?  (hh�e]r?  (hhe]r?  (jI>  ]r?  (h	h�e]r?  (hh�eeee]r?  (hheeej?  j?  ]r?  (j�,  ]r ?  (j�,  ]r!?  (j�,  ]r"?  (h	j�  e]r#?  (hh�e]r$?  (hhe]r%?  (jD>  ]r&?  (h	he]r'?  (hh�e]r(?  (hhe]r)?  (jI>  ]r*?  (h	h�e]r+?  (hh�eeee]r,?  (hheeej?  j?  j?  j?  ]r-?  (j�,  ]r.?  (j�,  ]r/?  (j�,  ]r0?  (h	j�  e]r1?  (hh�e]r2?  (hhe]r3?  (jD>  ]r4?  (h	he]r5?  (hh�e]r6?  (hhe]r7?  (jI>  ]r8?  (h	h�e]r9?  (hh�eeee]r:?  (hheeej-?  j-?  ]r;?  (j�,  ]r<?  (j�,  ]r=?  (j�,  ]r>?  (h	j�  e]r??  (hh�e]r@?  (hhe]rA?  (jD>  ]rB?  (h	he]rC?  (hh�e]rD?  (hhe]rE?  (jI>  ]rF?  (h	h�e]rG?  (hh�eeee]rH?  (hheee]rI?  (j�,  ]rJ?  (j�,  ]rK?  (j�,  ]rL?  (h	j�  e]rM?  (hh�e]rN?  (hhe]rO?  (jD>  ]rP?  (h	he]rQ?  (hh�e]rR?  (hhe]rS?  (jI>  ]rT?  (h	h�e]rU?  (hh�eeee]rV?  (hheee]rW?  (j�,  ]rX?  (j�,  ]rY?  (j�,  ]rZ?  (h	j�  e]r[?  (hh�e]r\?  (hhe]r]?  (jD>  ]r^?  (h	he]r_?  (hh�e]r`?  (hhe]ra?  (jI>  ]rb?  (h	h�e]rc?  (hh�eeee]rd?  (hheee]re?  (j�,  ]rf?  (j�,  ]rg?  (j�,  ]rh?  (h	j�  e]ri?  (hh�e]rj?  (hhe]rk?  (jD>  ]rl?  (h	he]rm?  (hh�e]rn?  (hhe]ro?  (jI>  ]rp?  (h	h�e]rq?  (hh�eeee]rr?  (hheeeje?  ]rs?  (j�,  ]rt?  (j�,  ]ru?  (j�,  ]rv?  (h	j�  e]rw?  (hh�e]rx?  (hhe]ry?  (jD>  ]rz?  (h	he]r{?  (hh�e]r|?  (hhe]r}?  (jI>  ]r~?  (h	h�e]r?  (hh�eeee]r�?  (hheeejs?  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (h	j�  e]r�?  (hh�e]r�?  (hhe]r�?  (jD>  ]r�?  (h	he]r�?  (hh�e]r�?  (hhe]r�?  (jI>  ]r�?  (h	h�e]r�?  (hh�eeee]r�?  (hheee]r�?  (j�,  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (h	j�  e]r�?  (hh�e]r�?  (hhe]r�?  (jD>  ]r�?  (h	he]r�?  (hh�e]r�?  (hhe]r�?  (jI>  ]r�?  (h	h�e]r�?  (hh�eeee]r�?  (hheeej�?  j�?  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (h	h�e]r�?  (hh�e]r�?  (hhe]r�?  (jD>  ]r�?  (h	he]r�?  (hh�e]r�?  (hhe]r�?  (jI>  ]r�?  (h	h�e]r�?  (hh�eeee]r�?  (hheeej�?  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (h	h�e]r�?  (hh�e]r�?  (hhe]r�?  (jD>  ]r�?  (h	he]r�?  (hh�e]r�?  (hhe]r�?  (jI>  ]r�?  (h	h�e]r�?  (hh�eeee]r�?  (hheee]r�?  (j�,  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (h	h�e]r�?  (hh�e]r�?  (hhe]r�?  (jD>  ]r�?  (h	he]r�?  (hh�e]r�?  (hhe]r�?  (jI>  ]r�?  (h	h�e]r�?  (hh�eeee]r�?  (hheeej�?  j�?  j�?  j�?  j�?  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (h	h�e]r�?  (hh�e]r�?  (hhe]r�?  (jD>  ]r�?  (h	he]r�?  (hh�e]r�?  (hhe]r�?  (jI>  ]r�?  (h	h�e]r�?  (hh�eeee]r�?  (hheeej�?  j�?  j�?  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (h	h�e]r�?  (hh�e]r�?  (hhe]r�?  (jD>  ]r�?  (h	he]r�?  (hh�e]r�?  (hhe]r�?  (jI>  ]r�?  (h	h�e]r�?  (hh�eeee]r�?  (hheeej�?  j�?  j�?  j�?  j�?  j�?  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (h	h�e]r�?  (hh�e]r�?  (hhe]r�?  (jD>  ]r�?  (h	he]r�?  (hh�e]r�?  (hhe]r�?  (jI>  ]r�?  (h	h�e]r�?  (hh�eeee]r�?  (hheee]r�?  (j�,  ]r�?  (j�,  ]r�?  (j�,  ]r�?  (h	h�e]r�?  (hh�e]r�?  (hhe]r�?  (jD>  ]r�?  (h	he]r�?  (hh�e]r�?  (hhe]r�?  (jI>  ]r�?  (h	h�e]r�?  (hh�eeee]r�?  (hheee]r�?  (j�,  ]r @  (j�,  ]r@  (j�,  ]r@  (h	h�e]r@  (hh�e]r@  (hhe]r@  (jD>  ]r@  (h	he]r@  (hh�e]r@  (hhe]r	@  (jI>  ]r
@  (h	h�e]r@  (hh�eeee]r@  (hheeej�?  j�?  j�?  j�?  j�?  j�?  j�?  j�?  j�?  j�?  j�?  ]r@  (j�,  ]r@  (j�,  ]r@  (j�,  ]r@  (h	j�  e]r@  (hh�e]r@  (hhe]r@  (jD>  ]r@  (h	he]r@  (hh�e]r@  (hhe]r@  (jI>  ]r@  (h	h�e]r@  (hh�eeee]r@  (hheeej@  j@  j@  j@  j@  ]r@  (j�,  ]r@  (j�,  ]r@  (j�,  ]r@  (h	h�e]r@  (hh�e]r @  (hhe]r!@  (jD>  ]r"@  (h	he]r#@  (hh�e]r$@  (hhe]r%@  (jI>  ]r&@  (h	h�e]r'@  (hh�eeee]r(@  (hheeej@  j@  j@  ]r)@  (j�,  ]r*@  (j�,  ]r+@  (j�,  ]r,@  (h	h�e]r-@  (hh�e]r.@  (hhe]r/@  (jD>  ]r0@  (h	he]r1@  (hh�e]r2@  (hhe]r3@  (jI>  ]r4@  (h	h�e]r5@  (hh�eeee]r6@  (hheeej)@  ]r7@  (j�,  ]r8@  (j�,  ]r9@  (j�,  ]r:@  (h	h�e]r;@  (hh�e]r<@  (hhe]r=@  (jD>  ]r>@  (h	he]r?@  (hh�e]r@@  (hhe]rA@  (jI>  ]rB@  (h	h�e]rC@  (hh�eeee]rD@  (hheeej7@  j7@  j7@  j7@  j7@  j7@  ]rE@  (j�,  ]rF@  (j�,  ]rG@  (j�,  ]rH@  (h	h�e]rI@  (hh�e]rJ@  (hhe]rK@  (jD>  ]rL@  (h	he]rM@  (hh�e]rN@  (hhe]rO@  (jI>  ]rP@  (h	h�e]rQ@  (hh�eeee]rR@  (hheeejE@  ]rS@  (j�,  ]rT@  (j�,  ]rU@  (j�,  ]rV@  (h	h�e]rW@  (hh�e]rX@  (hhe]rY@  (jD>  ]rZ@  (h	he]r[@  (hh�e]r\@  (hhe]r]@  (jI>  ]r^@  (h	h�e]r_@  (hh�eeee]r`@  (hheeejS@  jS@  jS@  jS@  jS@  jS@  jS@  jS@  jS@  jS@  jS@  jS@  jS@  jS@  jS@  jS@  ]ra@  (j�,  ]rb@  (j�,  ]rc@  (j�,  ]rd@  (h	h�e]re@  (hh�e]rf@  (hhe]rg@  (jD>  ]rh@  (h	he]ri@  (hh�e]rj@  (hhe]rk@  (jI>  ]rl@  (h	h�e]rm@  (hh�eeee]rn@  (hheee]ro@  (j�,  ]rp@  (j�,  ]rq@  (j�,  ]rr@  (h	h�e]rs@  (hh�e]rt@  (hhe]ru@  (jD>  ]rv@  (h	he]rw@  (hh�e]rx@  (hhe]ry@  (jI>  ]rz@  (h	h�e]r{@  (hh�eeee]r|@  (hheee]r}@  (j�,  ]r~@  (j�,  ]r@  (j�,  ]r�@  (h	h�e]r�@  (hh�e]r�@  (hhe]r�@  (jD>  ]r�@  (h	he]r�@  (hh�e]r�@  (hhe]r�@  (jI>  ]r�@  (h	h�e]r�@  (hh�eeee]r�@  (hheee]r�@  (j�,  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (h	h�e]r�@  (hh�e]r�@  (hhe]r�@  (jD>  ]r�@  (h	he]r�@  (hh�e]r�@  (hhe]r�@  (jI>  ]r�@  (h	h�e]r�@  (hh�eeee]r�@  (hheeej�@  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (h	h�e]r�@  (hh�e]r�@  (hhe]r�@  (jD>  ]r�@  (h	he]r�@  (hh�e]r�@  (hhe]r�@  (jI>  ]r�@  (h	h�e]r�@  (hh�eeee]r�@  (hheee]r�@  (j�,  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (h	h�e]r�@  (hh�e]r�@  (hhe]r�@  (jD>  ]r�@  (h	he]r�@  (hh�e]r�@  (hhe]r�@  (jI>  ]r�@  (h	h�e]r�@  (hh�eeee]r�@  (hheeej�@  j�@  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (h	h�e]r�@  (hh�e]r�@  (hhe]r�@  (jD>  ]r�@  (h	he]r�@  (hh�e]r�@  (hhe]r�@  (jI>  ]r�@  (h	h�e]r�@  (hh�eeee]r�@  (hheeej�@  j�@  j�@  j�@  j�@  j�@  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (h	h�e]r�@  (hh�e]r�@  (hhe]r�@  (jD>  ]r�@  (h	he]r�@  (hh�e]r�@  (hhe]r�@  (jI>  ]r�@  (h	h�e]r�@  (hh�eeee]r�@  (hheeej�@  j�@  j�@  j�@  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (h	h�e]r�@  (hh�e]r�@  (hhe]r�@  (jD>  ]r�@  (h	he]r�@  (hh�e]r�@  (hhe]r�@  (jI>  ]r�@  (h	h�e]r�@  (hh�eeee]r�@  (hheeej�@  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (h	h�e]r�@  (hh�e]r�@  (hhe]r�@  (jD>  ]r�@  (h	he]r�@  (hh�e]r�@  (hhe]r�@  (jI>  ]r�@  (h	h�e]r�@  (hh�eeee]r�@  (hheeej�@  j�@  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (h	h�e]r�@  (hh�e]r�@  (hhe]r�@  (jD>  ]r�@  (h	he]r�@  (hh�e]r�@  (hhe]r�@  (jI>  ]r�@  (h	h�e]r�@  (hh�eeee]r�@  (hheeej�@  j�@  j�@  j�@  j�@  j�@  j�@  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (j�,  ]r�@  (h	h�e]r�@  (hh�e]r A  (hhe]rA  (jD>  ]rA  (h	he]rA  (hh�e]rA  (hhe]rA  (jI>  ]rA  (h	h�e]rA  (hh�eeee]rA  (hheeej�@  j�@  j�@  j�@  ]r	A  (j�,  ]r
A  (j�,  ]rA  (j�,  ]rA  (h	j�  e]rA  (hh�e]rA  (hhe]rA  (jD>  ]rA  (h	he]rA  (hh�e]rA  (hhe]rA  (jI>  ]rA  (h	h�e]rA  (hh�eeee]rA  (hheeej	A  j	A  j	A  j	A  ]rA  (j�,  ]rA  (j�,  ]rA  (j�,  ]rA  (h	j�  e]rA  (hh�e]rA  (hhe]rA  (jD>  ]rA  (h	he]rA  (hh�e]r A  (hhe]r!A  (jI>  ]r"A  (h	h�e]r#A  (hh�eeee]r$A  (hheeejA  jA  ]r%A  (j�,  ]r&A  (j�,  ]r'A  (j�,  ]r(A  (h	h�e]r)A  (hh�e]r*A  (hhe]r+A  (jD>  ]r,A  (h	he]r-A  (hh�e]r.A  (hhe]r/A  (jI>  ]r0A  (h	h�e]r1A  (hh�eeee]r2A  (hheeej%A  j%A  ]r3A  (j�,  ]r4A  (j�,  ]r5A  (j�,  ]r6A  (h	h�e]r7A  (hh�e]r8A  (hhe]r9A  (jD>  ]r:A  (h	he]r;A  (hh�e]r<A  (hhe]r=A  (jI>  ]r>A  (h	h�e]r?A  (hh�eeee]r@A  (hheeej3A  ]rAA  (j�,  ]rBA  (j�,  ]rCA  (j�,  ]rDA  (h	j�  e]rEA  (hh�e]rFA  (hhe]rGA  (jD>  ]rHA  (h	he]rIA  (hh�e]rJA  (hhe]rKA  (jI>  ]rLA  (h	h�e]rMA  (hh�eeee]rNA  (hheeejAA  jAA  ]rOA  (j�,  ]rPA  (j�,  ]rQA  (j�,  ]rRA  (h	j�  e]rSA  (hh�e]rTA  (hhe]rUA  (jD>  ]rVA  (h	he]rWA  (hh�e]rXA  (hhe]rYA  (jI>  ]rZA  (h	h�e]r[A  (hh�eeee]r\A  (hheeejOA  jOA  ]r]A  (j�,  ]r^A  (j�,  ]r_A  (j�,  ]r`A  (h	j�  e]raA  (hh�e]rbA  (hhe]rcA  (jD>  ]rdA  (h	he]reA  (hh�e]rfA  (hhe]rgA  (jI>  ]rhA  (h	h�e]riA  (hh�eeee]rjA  (hheeej]A  j]A  j]A  j]A  j]A  j]A  j]A  j]A  j]A  j]A  j]A  j]A  j]A  j]A  j]A  ]rkA  (j�,  ]rlA  (j�,  ]rmA  (j�,  ]rnA  (h	j�  e]roA  (hh�e]rpA  (hhe]rqA  (jD>  ]rrA  (h	he]rsA  (hh�e]rtA  (hhe]ruA  (jI>  ]rvA  (h	h�e]rwA  (hh�eeee]rxA  (hheeejkA  jkA  jkA  jkA  ]ryA  (j�,  ]rzA  (j�,  ]r{A  (j�,  ]r|A  (h	j�  e]r}A  (hh�e]r~A  (hhe]rA  (jD>  ]r�A  (h	he]r�A  (hh�e]r�A  (hhe]r�A  (jI>  ]r�A  (h	h�e]r�A  (hh�eeee]r�A  (hheee]r�A  (j�,  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (h	h�e]r�A  (hh�e]r�A  (hhe]r�A  (jD>  ]r�A  (h	he]r�A  (hh�e]r�A  (hhe]r�A  (jI>  ]r�A  (h	h�e]r�A  (hh�eeee]r�A  (hheeej�A  j�A  j�A  j�A  j�A  j�A  j�A  j�A  j�A  j�A  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (h	h�e]r�A  (hh�e]r�A  (hhe]r�A  (jD>  ]r�A  (h	he]r�A  (hh�e]r�A  (hhe]r�A  (jI>  ]r�A  (h	h�e]r�A  (hh�eeee]r�A  (hheee]r�A  (j�,  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (h	h�e]r�A  (hh�e]r�A  (hhe]r�A  (jD>  ]r�A  (h	he]r�A  (hh�e]r�A  (hhe]r�A  (jI>  ]r�A  (h	h�e]r�A  (hh�eeee]r�A  (hheeej�A  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (h	h�e]r�A  (hh�e]r�A  (hhe]r�A  (jD>  ]r�A  (h	he]r�A  (hh�e]r�A  (hhe]r�A  (jI>  ]r�A  (h	h�e]r�A  (hh�eeee]r�A  (hheeej�A  j�A  j�A  j�A  j�A  j�A  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (h	h�e]r�A  (hh�e]r�A  (hhe]r�A  (jD>  ]r�A  (h	he]r�A  (hh�e]r�A  (hhe]r�A  (jI>  ]r�A  (h	h�e]r�A  (hh�eeee]r�A  (hheeej�A  j�A  j�A  j�A  j�A  j�A  j�A  j�A  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (h	h�e]r�A  (hh�e]r�A  (hhe]r�A  (jD>  ]r�A  (h	he]r�A  (hh�e]r�A  (hhe]r�A  (jI>  ]r�A  (h	h�e]r�A  (hh�eeee]r�A  (hheeej�A  j�A  j�A  j�A  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (h	h�e]r�A  (hh�e]r�A  (hhe]r�A  (jD>  ]r�A  (h	he]r�A  (hh�e]r�A  (hhe]r�A  (jI>  ]r�A  (h	h�e]r�A  (hh�eeee]r�A  (hheee]r�A  (j�,  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (h	h�e]r�A  (hh�e]r�A  (hhe]r�A  (jD>  ]r�A  (h	he]r�A  (hh�e]r�A  (hhe]r�A  (jI>  ]r�A  (h	h�e]r�A  (hh�eeee]r�A  (hheee]r�A  (j�,  ]r�A  (j�,  ]r�A  (j�,  ]r�A  (h	h�e]r�A  (hh�e]r�A  (hhe]r�A  (jD>  ]r�A  (h	he]r�A  (hh�e]r B  (hhe]rB  (jI>  ]rB  (h	h�e]rB  (hh�eeee]rB  (hheeej�A  ]rB  (j�,  ]rB  (j�,  ]rB  (j�,  ]rB  (h	h�e]r	B  (hh�e]r
B  (hhe]rB  (jD>  ]rB  (h	he]rB  (hh�e]rB  (hhe]rB  (jI>  ]rB  (h	h�e]rB  (hh�eeee]rB  (hheeejB  jB  jB  jB  ]rB  (j�,  ]rB  (j�,  ]rB  (j�,  ]rB  (h	h�e]rB  (hh�e]rB  (hhe]rB  (jD>  ]rB  (h	he]rB  (hh�e]rB  (hhe]rB  (jI>  ]rB  (h	h�e]rB  (hh�eeee]r B  (hheeejB  jB  jB  ]r!B  (j�,  ]r"B  (j�,  ]r#B  (j�,  ]r$B  (h	h�e]r%B  (hh�e]r&B  (hhe]r'B  (jD>  ]r(B  (h	he]r)B  (hh�e]r*B  (hhe]r+B  (jI>  ]r,B  (h	h�e]r-B  (hh�eeee]r.B  (hheeej!B  j!B  j!B  j!B  ]r/B  (j�,  ]r0B  (j�,  ]r1B  (j�,  ]r2B  (h	h�e]r3B  (hh�e]r4B  (hhe]r5B  (jD>  ]r6B  (h	he]r7B  (hh�e]r8B  (hhe]r9B  (jI>  ]r:B  (h	h�e]r;B  (hh�eeee]r<B  (hheeej/B  j/B  j/B  ]r=B  (j�,  ]r>B  (j�,  ]r?B  (j�,  ]r@B  (h	h�e]rAB  (hh�e]rBB  (hhe]rCB  (jD>  ]rDB  (h	he]rEB  (hh�e]rFB  (hhe]rGB  (jI>  ]rHB  (h	h�e]rIB  (hh�eeee]rJB  (hheeej=B  j=B  j=B  j=B  j=B  j=B  j=B  ]rKB  (j�,  ]rLB  (j�,  ]rMB  (j�,  ]rNB  (h	h�e]rOB  (hh�e]rPB  (hhe]rQB  (jD>  ]rRB  (h	he]rSB  (hh�e]rTB  (hhe]rUB  (jI>  ]rVB  (h	h�e]rWB  (hh�eeee]rXB  (hheeejKB  jKB  jKB  jKB  jKB  ]rYB  (j�,  ]rZB  (j�,  ]r[B  (j�,  ]r\B  (h	h�e]r]B  (hh�e]r^B  (hhe]r_B  (jD>  ]r`B  (h	he]raB  (hh�e]rbB  (hhe]rcB  (jI>  ]rdB  (h	h�e]reB  (hh�eeee]rfB  (hheeejYB  jYB  ]rgB  (j�,  ]rhB  (j�,  ]riB  (j�,  ]rjB  (h	h�e]rkB  (hh�e]rlB  (hhe]rmB  (jD>  ]rnB  (h	he]roB  (hh�e]rpB  (hhe]rqB  (jI>  ]rrB  (h	h�e]rsB  (hh�eeee]rtB  (hheeejgB  jgB  jgB  ]ruB  (j�,  ]rvB  (j�,  ]rwB  (j�,  ]rxB  (h	h�e]ryB  (hh�e]rzB  (hhe]r{B  (jD>  ]r|B  (h	he]r}B  (hh�e]r~B  (hhe]rB  (jI>  ]r�B  (h	h�e]r�B  (hh�eeee]r�B  (hheeejuB  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (h	h�e]r�B  (hh�e]r�B  (hhe]r�B  (jD>  ]r�B  (h	he]r�B  (hh�e]r�B  (hhe]r�B  (jI>  ]r�B  (h	h�e]r�B  (hh�eeee]r�B  (hheeej�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (h	h�e]r�B  (hh�e]r�B  (hhe]r�B  (jD>  ]r�B  (h	he]r�B  (hh�e]r�B  (hhe]r�B  (jI>  ]r�B  (h	h�e]r�B  (hh�eeee]r�B  (hheeej�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  j�B  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (h	h�e]r�B  (hh�e]r�B  (hhe]r�B  (jD>  ]r�B  (h	he]r�B  (hh�e]r�B  (hhe]r�B  (jI>  ]r�B  (h	h�e]r�B  (hh�eeee]r�B  (hheeej�B  j�B  j�B  j�B  j�B  j�B  j�B  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (h	h�e]r�B  (hh�e]r�B  (hhe]r�B  (jD>  ]r�B  (h	he]r�B  (hh�e]r�B  (hhe]r�B  (jI>  ]r�B  (h	h�e]r�B  (hh�eeee]r�B  (hheeej�B  j�B  j�B  j�B  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (h	h�e]r�B  (hh�e]r�B  (hhe]r�B  (jD>  ]r�B  (h	he]r�B  (hh�e]r�B  (hhe]r�B  (jI>  ]r�B  (h	h�e]r�B  (hh�eeee]r�B  (hheeej�B  j�B  j�B  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (h	h�e]r�B  (hh�e]r�B  (hhe]r�B  (jD>  ]r�B  (h	he]r�B  (hh�e]r�B  (hhe]r�B  (jI>  ]r�B  (h	h�e]r�B  (hh�eeee]r�B  (hheeej�B  j�B  j�B  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (h	h�e]r�B  (hh�e]r�B  (hhe]r�B  (jD>  ]r�B  (h	he]r�B  (hh�e]r�B  (hhe]r�B  (jI>  ]r�B  (h	h�e]r�B  (hh�eeee]r�B  (hheeej�B  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (h	h�e]r�B  (hh�e]r�B  (hhe]r�B  (jD>  ]r�B  (h	he]r�B  (hh�e]r�B  (hhe]r�B  (jI>  ]r�B  (h	h�e]r�B  (hh�eeee]r�B  (hheeej�B  j�B  j�B  j�B  j�B  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (j�,  ]r�B  (h	h�e]r�B  (hh�e]r�B  (hhe]r�B  (jD>  ]r�B  (h	he]r�B  (hh�e]r�B  (hhe]r�B  (jI>  ]r�B  (h	h�e]r�B  (hh�eeee]r C  (hheeej�B  j�B  j�B  j�B  j�B  j�B  ]rC  (j�,  ]rC  (j�,  ]rC  (j�,  ]rC  (h	h�e]rC  (hh�e]rC  (hhe]rC  (jD>  ]rC  (h	he]r	C  (hh�e]r
C  (hhe]rC  (jI>  ]rC  (h	h�e]rC  (hh�eeee]rC  (hheeejC  jC  jC  jC  jC  jC  ]rC  (j�,  ]rC  (j�,  ]rC  (j�,  ]rC  (h	h�e]rC  (hh�e]rC  (hhe]rC  (jD>  ]rC  (h	he]rC  (hh�e]rC  (hhe]rC  (jI>  ]rC  (h	h�e]rC  (hh�eeee]rC  (hheeejC  ]rC  (j�,  ]rC  (j�,  ]rC  (j�,  ]r C  (h	h�e]r!C  (hh�e]r"C  (hhe]r#C  (jD>  ]r$C  (h	he]r%C  (hh�e]r&C  (hhe]r'C  (jI>  ]r(C  (h	h�e]r)C  (hh�eeee]r*C  (hheeejC  ]r+C  (j�,  ]r,C  (j�,  ]r-C  (j�,  ]r.C  (h	h�e]r/C  (hh�e]r0C  (hhe]r1C  (jD>  ]r2C  (h	he]r3C  (hh�e]r4C  (hhe]r5C  (jI>  ]r6C  (h	h�e]r7C  (hh�eeee]r8C  (hheeej+C  j+C  j+C  ]r9C  (j�,  ]r:C  (j�,  ]r;C  (j�,  ]r<C  (h	h�e]r=C  (hh�e]r>C  (hhe]r?C  (jD>  ]r@C  (h	he]rAC  (hh�e]rBC  (hhe]rCC  (jI>  ]rDC  (h	h�e]rEC  (hh�eeee]rFC  (hheeej9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  j9C  ]rGC  (j�,  ]rHC  (j�,  ]rIC  (j�,  ]rJC  (h	h�e]rKC  (hh�e]rLC  (hhe]rMC  (jD>  ]rNC  (h	he]rOC  (hh�e]rPC  (hhe]rQC  (jI>  ]rRC  (h	h�e]rSC  (hh�eeee]rTC  (hheeejGC  jGC  jGC  jGC  jGC  ]rUC  (j�,  ]rVC  (j�,  ]rWC  (j�,  ]rXC  (h	h�e]rYC  (hh�e]rZC  (hhe]r[C  (jD>  ]r\C  (h	he]r]C  (hh�e]r^C  (hhe]r_C  (jI>  ]r`C  (h	h�e]raC  (hh�eeee]rbC  (hheeejUC  jUC  ]rcC  (j�,  ]rdC  (j�,  ]reC  (j�,  ]rfC  (h	h�e]rgC  (hh�e]rhC  (hhe]riC  (jD>  ]rjC  (h	he]rkC  (hh�e]rlC  (hhe]rmC  (jI>  ]rnC  (h	h�e]roC  (hh�eeee]rpC  (hheeejcC  ]rqC  (j�,  ]rrC  (j�,  ]rsC  (j�,  ]rtC  (h	h�e]ruC  (hh�e]rvC  (hhe]rwC  (jD>  ]rxC  (h	he]ryC  (hh�e]rzC  (hhe]r{C  (jI>  ]r|C  (h	h�e]r}C  (hh�eeee]r~C  (hheeejqC  jqC  jqC  jqC  jqC  jqC  jqC  jqC  jqC  jqC  jqC  jqC  jqC  jqC  jqC  jqC  ]rC  (j�,  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (h	h�e]r�C  (hh�e]r�C  (hhe]r�C  (jD>  ]r�C  (h	he]r�C  (hh�e]r�C  (hhe]r�C  (jI>  ]r�C  (h	h�e]r�C  (hh�eeee]r�C  (hheeejC  jC  jC  jC  jC  jC  jC  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (h	h�e]r�C  (hh�e]r�C  (hhe]r�C  (jD>  ]r�C  (h	he]r�C  (hh�e]r�C  (hhe]r�C  (jI>  ]r�C  (h	h�e]r�C  (hh�eeee]r�C  (hheeej�C  j�C  j�C  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (h	h�e]r�C  (hh�e]r�C  (hhe]r�C  (jD>  ]r�C  (h	he]r�C  (hh�e]r�C  (hhe]r�C  (jI>  ]r�C  (h	h�e]r�C  (hh�eeee]r�C  (hheeej�C  j�C  j�C  j�C  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (h	h�e]r�C  (hh�e]r�C  (hhe]r�C  (jD>  ]r�C  (h	he]r�C  (hh�e]r�C  (hhe]r�C  (jI>  ]r�C  (h	h�e]r�C  (hh�eeee]r�C  (hheeej�C  j�C  j�C  j�C  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (h	h�e]r�C  (hh�e]r�C  (hhe]r�C  (jD>  ]r�C  (h	he]r�C  (hh�e]r�C  (hhe]r�C  (jI>  ]r�C  (h	h�e]r�C  (hh�eeee]r�C  (hheee]r�C  (j�,  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (h	h�e]r�C  (hh�e]r�C  (hhe]r�C  (jD>  ]r�C  (h	he]r�C  (hh�e]r�C  (hhe]r�C  (jI>  ]r�C  (h	h�e]r�C  (hh�eeee]r�C  (hheeej�C  j�C  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (h	j�  e]r�C  (hh�e]r�C  (hhe]r�C  (jD>  ]r�C  (h	he]r�C  (hh�e]r�C  (hhe]r�C  (jI>  ]r�C  (h	h�e]r�C  (hh�eeee]r�C  (hheeej�C  j�C  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (h	j�  e]r�C  (hh�e]r�C  (hhe]r�C  (jD>  ]r�C  (h	he]r�C  (hh�e]r�C  (hhe]r�C  (jI>  ]r�C  (h	h�e]r�C  (hh�eeee]r�C  (hheeej�C  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (h	j�  e]r�C  (hh�e]r�C  (hhe]r�C  (jD>  ]r�C  (h	he]r�C  (hh�e]r�C  (hhe]r�C  (jI>  ]r�C  (h	h�e]r�C  (hh�eeee]r�C  (hheeej�C  j�C  ]r�C  (j�,  ]r�C  (j�,  ]r�C  (j�,  ]r D  (h	j�  e]rD  (hh�e]rD  (hhe]rD  (jD>  ]rD  (h	he]rD  (hh�e]rD  (hhe]rD  (jI>  ]rD  (h	h�e]r	D  (hh�eeee]r
D  (hheee]rD  (j�,  ]rD  (j�,  ]rD  (j�,  ]rD  (h	j�  e]rD  (hh�e]rD  (hhe]rD  (jD>  ]rD  (h	he]rD  (hh�e]rD  (hhe]rD  (jI>  ]rD  (h	h�e]rD  (hh�eeee]rD  (hheeejD  jD  ]rD  (j�,  ]rD  (j�,  ]rD  (j�,  ]rD  (h	h�e]rD  (hh�e]rD  (hhe]rD  (jD>  ]r D  (h	he]r!D  (hh�e]r"D  (hhe]r#D  (jI>  ]r$D  (h	h�e]r%D  (hh�eeee]r&D  (hheee]r'D  (j�,  ]r(D  (j�,  ]r)D  (j�,  ]r*D  (h	h�e]r+D  (hh�e]r,D  (hhe]r-D  (jD>  ]r.D  (h	he]r/D  (hh�e]r0D  (hhe]r1D  (jI>  ]r2D  (h	h�e]r3D  (hh�eeee]r4D  (hheeej'D  j'D  j'D  j'D  ]r5D  (j�,  ]r6D  (j�,  ]r7D  (j�,  ]r8D  (h	h�e]r9D  (hh�e]r:D  (hhe]r;D  (jD>  ]r<D  (h	he]r=D  (hh�e]r>D  (hhe]r?D  (jI>  ]r@D  (h	h�e]rAD  (hh�eeee]rBD  (hheeej5D  ]rCD  (j�,  ]rDD  (j�,  ]rED  (j�,  ]rFD  (h	h�e]rGD  (hh�e]rHD  (hhe]rID  (jD>  ]rJD  (h	he]rKD  (hh�e]rLD  (hhe]rMD  (jI>  ]rND  (h	h�e]rOD  (hh�eeee]rPD  (hheeejCD  ]rQD  (j�,  ]rRD  (j�,  ]rSD  (j�,  ]rTD  (h	h�e]rUD  (hh�e]rVD  (hhe]rWD  (jD>  ]rXD  (h	he]rYD  (hh�e]rZD  (hhe]r[D  (jI>  ]r\D  (h	h�e]r]D  (hh�eeee]r^D  (hheeejQD  jQD  jQD  jQD  jQD  jQD  ]r_D  (j�,  ]r`D  (j�,  ]raD  (j�,  ]rbD  (h	h�e]rcD  (hh�e]rdD  (hhe]reD  (jD>  ]rfD  (h	he]rgD  (hh�e]rhD  (hhe]riD  (jI>  ]rjD  (h	h�e]rkD  (hh�eeee]rlD  (hheeej_D  j_D  j_D  j_D  j_D  j_D  ]rmD  (j�,  ]rnD  (j�,  ]roD  (j�,  ]rpD  (h	h�e]rqD  (hh�e]rrD  (hhe]rsD  (jD>  ]rtD  (h	he]ruD  (hh�e]rvD  (hhe]rwD  (jI>  ]rxD  (h	h�e]ryD  (hh�eeee]rzD  (hheeejmD  ]r{D  (j�,  ]r|D  (j�,  ]r}D  (j�,  ]r~D  (h	h�e]rD  (hh�e]r�D  (hhe]r�D  (jD>  ]r�D  (h	he]r�D  (hh�e]r�D  (hhe]r�D  (jI>  ]r�D  (h	h�e]r�D  (hh�eeee]r�D  (hheeej{D  j{D  j{D  j{D  j{D  j{D  j{D  j{D  j{D  j{D  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (h	h�e]r�D  (hh�e]r�D  (hhe]r�D  (jD>  ]r�D  (h	he]r�D  (hh�e]r�D  (hhe]r�D  (jI>  ]r�D  (h	h�e]r�D  (hh�eeee]r�D  (hheee]r�D  (j�,  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (h	h�e]r�D  (hh�e]r�D  (hhe]r�D  (jD>  ]r�D  (h	he]r�D  (hh�e]r�D  (hhe]r�D  (jI>  ]r�D  (h	h�e]r�D  (hh�eeee]r�D  (hheeej�D  j�D  j�D  j�D  j�D  j�D  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (h	h�e]r�D  (hh�e]r�D  (hhe]r�D  (jD>  ]r�D  (h	he]r�D  (hh�e]r�D  (hhe]r�D  (jI>  ]r�D  (h	h�e]r�D  (hh�eeee]r�D  (hheee]r�D  (j�,  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (h	h�e]r�D  (hh�e]r�D  (hhe]r�D  (jD>  ]r�D  (h	he]r�D  (hh�e]r�D  (hhe]r�D  (jI>  ]r�D  (h	h�e]r�D  (hh�eeee]r�D  (hheee]r�D  (j�,  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (h	h�e]r�D  (hh�e]r�D  (hhe]r�D  (jD>  ]r�D  (h	he]r�D  (hh�e]r�D  (hhe]r�D  (jI>  ]r�D  (h	h�e]r�D  (hh�eeee]r�D  (hheeej�D  j�D  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (h	j�  e]r�D  (hh�e]r�D  (hhe]r�D  (jD>  ]r�D  (h	he]r�D  (hh�e]r�D  (hhe]r�D  (jI>  ]r�D  (h	h�e]r�D  (hh�eeee]r�D  (hheeej�D  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (h	j�  e]r�D  (hh�e]r�D  (hhe]r�D  (jD>  ]r�D  (h	he]r�D  (hh�e]r�D  (hhe]r�D  (jI>  ]r�D  (h	h�e]r�D  (hh�eeee]r�D  (hheeej�D  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (h	j�  e]r�D  (hh�e]r�D  (hhe]r�D  (jD>  ]r�D  (h	he]r�D  (hh�e]r�D  (hhe]r�D  (jI>  ]r�D  (h	h�e]r�D  (hh�eeee]r�D  (hheeej�D  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (j�,  ]r�D  (h	j�  e]r�D  (hh�e]r�D  (hhe]r�D  (jD>  ]r E  (h	he]rE  (hh�e]rE  (hhe]rE  (jI>  ]rE  (h	h�e]rE  (hh�eeee]rE  (hheee]rE  (j�,  ]rE  (j�,  ]r	E  (j�,  ]r
E  (h	j�  e]rE  (hh�e]rE  (hhe]rE  (jD>  ]rE  (h	he]rE  (hh�e]rE  (hhe]rE  (jI>  ]rE  (h	h�e]rE  (hh�eeee]rE  (hheeejE  jE  jE  ]rE  (j�,  ]rE  (j�,  ]rE  (j�,  ]rE  (h	h�e]rE  (hh�e]rE  (hhe]rE  (jD>  ]rE  (h	he]rE  (hh�e]rE  (hhe]rE  (jI>  ]r E  (h	h�e]r!E  (hh�eeee]r"E  (hheeejE  jE  ]r#E  (j�,  ]r$E  (j�,  ]r%E  (j�,  ]r&E  (h	h�e]r'E  (hh�e]r(E  (hhe]r)E  (jD>  ]r*E  (h	he]r+E  (hh�e]r,E  (hhe]r-E  (jI>  ]r.E  (h	h�e]r/E  (hh�eeee]r0E  (hheee]r1E  (j�,  ]r2E  (j�,  ]r3E  (j�,  ]r4E  (h	h�e]r5E  (hh�e]r6E  (hhe]r7E  (jD>  ]r8E  (h	he]r9E  (hh�e]r:E  (hhe]r;E  (jI>  ]r<E  (h	h�e]r=E  (hh�eeee]r>E  (hheeej1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  j1E  ]r?E  (j�,  ]r@E  (j�,  ]rAE  (j�,  ]rBE  (h	h�e]rCE  (hh�e]rDE  (hhe]rEE  (jD>  ]rFE  (h	he]rGE  (hh�e]rHE  (hhe]rIE  (jI>  ]rJE  (h	h�e]rKE  (hh�eeee]rLE  (hheee]rME  (j�,  ]rNE  (j�,  ]rOE  (j�,  ]rPE  (h	h�e]rQE  (hh�e]rRE  (hhe]rSE  (jD>  ]rTE  (h	he]rUE  (hh�e]rVE  (hhe]rWE  (jI>  ]rXE  (h	h�e]rYE  (hh�eeee]rZE  (hheee]r[E  (j�,  ]r\E  (j�,  ]r]E  (j�,  ]r^E  (h	h�e]r_E  (hh�e]r`E  (hhe]raE  (jD>  ]rbE  (h	he]rcE  (hh�e]rdE  (hhe]reE  (jI>  ]rfE  (h	h�e]rgE  (hh�eeee]rhE  (hheeej[E  j[E  j[E  j[E  ]riE  (j�,  ]rjE  (j�,  ]rkE  (j�,  ]rlE  (h	h�e]rmE  (hh�e]rnE  (hhe]roE  (jD>  ]rpE  (h	he]rqE  (hh�e]rrE  (hhe]rsE  (jI>  ]rtE  (h	h�e]ruE  (hh�eeee]rvE  (hheeejiE  jiE  jiE  ]rwE  (j�,  ]rxE  (j�,  ]ryE  (j�,  ]rzE  (h	h�e]r{E  (hh�e]r|E  (hhe]r}E  (jD>  ]r~E  (h	he]rE  (hh�e]r�E  (hhe]r�E  (jI>  ]r�E  (h	h�e]r�E  (hh�eeee]r�E  (hheeejwE  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (h	h�e]r�E  (hh�e]r�E  (hhe]r�E  (jD>  ]r�E  (h	he]r�E  (hh�e]r�E  (hhe]r�E  (jI>  ]r�E  (h	h�e]r�E  (hh�eeee]r�E  (hheee]r�E  (j�,  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (h	h�e]r�E  (hh�e]r�E  (hhe]r�E  (jD>  ]r�E  (h	he]r�E  (hh�e]r�E  (hhe]r�E  (jI>  ]r�E  (h	h�e]r�E  (hh�eeee]r�E  (hheeej�E  j�E  j�E  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (h	j�  e]r�E  (hh�e]r�E  (hhe]r�E  (jD>  ]r�E  (h	he]r�E  (hh�e]r�E  (hhe]r�E  (jI>  ]r�E  (h	h�e]r�E  (hh�eeee]r�E  (hheeej�E  j�E  j�E  j�E  j�E  j�E  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (h	j�  e]r�E  (hh�e]r�E  (hhe]r�E  (jD>  ]r�E  (h	he]r�E  (hh�e]r�E  (hhe]r�E  (jI>  ]r�E  (h	h�e]r�E  (hh�eeee]r�E  (hheee]r�E  (j�,  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (h	j�  e]r�E  (hh�e]r�E  (hhe]r�E  (jD>  ]r�E  (h	he]r�E  (hh�e]r�E  (hhe]r�E  (jI>  ]r�E  (h	h�e]r�E  (hh�eeee]r�E  (hheeej�E  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (h	j�  e]r�E  (hh�e]r�E  (hhe]r�E  (jD>  ]r�E  (h	he]r�E  (hh�e]r�E  (hhe]r�E  (jI>  ]r�E  (h	h�e]r�E  (hh�eeee]r�E  (hheeej�E  j�E  j�E  j�E  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (h	j�  e]r�E  (hh�e]r�E  (hhe]r�E  (jD>  ]r�E  (h	he]r�E  (hh�e]r�E  (hhe]r�E  (jI>  ]r�E  (h	h�e]r�E  (hh�eeee]r�E  (hheeej�E  j�E  j�E  j�E  j�E  j�E  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (h	j�  e]r�E  (hh�e]r�E  (hhe]r�E  (jD>  ]r�E  (h	he]r�E  (hh�e]r�E  (hhe]r�E  (jI>  ]r�E  (h	h�e]r�E  (hh�eeee]r�E  (hheeej�E  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (j�,  ]r�E  (h	j�  e]r�E  (hh�e]r�E  (hhe]r�E  (jD>  ]r�E  (h	he]r�E  (hh�e]r�E  (hhe]r�E  (jI>  ]r F  (h	h�e]rF  (hh�eeee]rF  (hheeej�E  j�E  j�E  j�E  j�E  j�E  j�E  j�E  ]rF  (j�,  ]rF  (j�,  ]rF  (j�,  ]rF  (h	j�  e]rF  (hh�e]rF  (hhe]r	F  (jD>  ]r
F  (h	he]rF  (hh�e]rF  (hhe]rF  (jI>  ]rF  (h	h�e]rF  (hh�eeee]rF  (hheeejF  jF  jF  jF  jF  jF  jF  ]rF  (j�,  ]rF  (j�,  ]rF  (j�,  ]rF  (h	j�  e]rF  (hh�e]rF  (hhe]rF  (jD>  ]rF  (h	he]rF  (hh�e]rF  (hhe]rF  (jI>  ]rF  (h	h�e]rF  (hh�eeee]rF  (hheeejF  jF  jF  jF  jF  jF  jF  ]rF  (j�,  ]r F  (j�,  ]r!F  (j�,  ]r"F  (h	j�  e]r#F  (hh�e]r$F  (hhe]r%F  (jD>  ]r&F  (h	he]r'F  (hh�e]r(F  (hhe]r)F  (jI>  ]r*F  (h	h�e]r+F  (hh�eeee]r,F  (hheeejF  jF  jF  jF  jF  jF  ]r-F  (j�,  ]r.F  (j�,  ]r/F  (j�,  ]r0F  (h	j�  e]r1F  (hh�e]r2F  (hhe]r3F  (jD>  ]r4F  (h	he]r5F  (hh�e]r6F  (hhe]r7F  (jI>  ]r8F  (h	h�e]r9F  (hh�eeee]r:F  (hheee]r;F  (j�,  ]r<F  (j�,  ]r=F  (j�,  ]r>F  (h	j�  e]r?F  (hh�e]r@F  (hhe]rAF  (jD>  ]rBF  (h	he]rCF  (hh�e]rDF  (hhe]rEF  (jI>  ]rFF  (h	h�e]rGF  (hh�eeee]rHF  (hheeej;F  j;F  j;F  j;F  j;F  j;F  j;F  j;F  ]rIF  (j�,  ]rJF  (j�,  ]rKF  (j�,  ]rLF  (h	j�  e]rMF  (hh�e]rNF  (hhe]rOF  (jD>  ]rPF  (h	he]rQF  (hh�e]rRF  (hhe]rSF  (jI>  ]rTF  (h	h�e]rUF  (hh�eeee]rVF  (hheeejIF  jIF  e(jIF  e]rWF  (]rXF  (X   NormrYF  ]rZF  (X   Oblr[F  ]r\F  (X   Movedr]F  ]r^F  (h	X   anyr_F  e]r`F  (hX   squareraF  e]rbF  (hhe]rcF  (X   MovedrdF  ]reF  (h	he]rfF  (hX   anyrgF  e]rhF  (hhe]riF  (X	   Next-MoverjF  ]rkF  (h	X   anyrlF  e]rmF  (hX   squarernF  eeee]roF  (hheeejXF  ]rpF  (jYF  ]rqF  (j[F  ]rrF  (j]F  ]rsF  (h	j_F  e]rtF  (hjaF  e]ruF  (hhe]rvF  (jdF  ]rwF  (h	he]rxF  (hjgF  e]ryF  (hhe]rzF  (jjF  ]r{F  (h	jlF  e]r|F  (hh�eeee]r}F  (hheee]r~F  (jYF  ]rF  (j[F  ]r�F  (j]F  ]r�F  (h	j_F  e]r�F  (hjaF  e]r�F  (hhe]r�F  (jdF  ]r�F  (h	he]r�F  (hjgF  e]r�F  (hhe]r�F  (jjF  ]r�F  (h	jlF  e]r�F  (hh�eeee]r�F  (hheeej~F  j~F  j~F  j~F  j~F  j~F  j~F  ]r�F  (jYF  ]r�F  (j[F  ]r�F  (j]F  ]r�F  (h	j_F  e]r�F  (hjaF  e]r�F  (hhe]r�F  (jdF  ]r�F  (h	he]r�F  (hjgF  e]r�F  (hhe]r�F  (jjF  ]r�F  (h	jlF  e]r�F  (hh�eeee]r�F  (hheeej�F  ]r�F  (jYF  ]r�F  (j[F  ]r�F  (j]F  ]r�F  (h	j_F  e]r�F  (hh�e]r�F  (hhe]r�F  (jdF  ]r�F  (h	he]r�F  (hjgF  e]r�F  (hhe]r�F  (jjF  ]r�F  (h	jlF  e]r�F  (hh�eeee]r�F  (hheeej�F  j�F  j�F  ]r�F  (jYF  ]r�F  (j[F  ]r�F  (j]F  ]r�F  (h	j_F  e]r�F  (hh�e]r�F  (hhe]r�F  (jdF  ]r�F  (h	he]r�F  (hjgF  e]r�F  (hhe]r�F  (jjF  ]r�F  (h	jlF  e]r�F  (hh�eeee]r�F  (hheeej�F  j�F  j�F  j�F  j�F  j�F  ]r�F  (jYF  ]r�F  (j[F  ]r�F  (j]F  ]r�F  (h	j_F  e]r�F  (hh�e]r�F  (hhe]r�F  (jdF  ]r�F  (h	he]r�F  (hh�e]r�F  (hhe]r�F  (jjF  ]r�F  (h	jlF  e]r�F  (hh�eeee]r�F  (hheeej�F  ]r�F  (jYF  ]r�F  (j[F  ]r�F  (j]F  ]r�F  (h	j_F  e]r�F  (hh�e]r�F  (hhe]r�F  (jdF  ]r�F  (h	he]r�F  (hh�e]r�F  (hhe]r�F  (jjF  ]r�F  (h	jlF  e]r�F  (hh�eeee]r�F  (hheeej�F  ]r�F  (jYF  ]r�F  (j[F  ]r�F  (j]F  ]r�F  (h	j_F  e]r�F  (hh�e]r�F  (hhe]r�F  (jdF  ]r�F  (h	he]r�F  (hh�e]r�F  (hhe]r�F  (jjF  ]r�F  (h	jlF  e]r�F  (hh�eeee]r�F  (hheeej�F  j�F  j�F  j�F  j�F  j�F  j�F  ]r�F  (jYF  ]r�F  (j[F  ]r�F  (j]F  ]r�F  (h	j_F  e]r�F  (hh�e]r�F  (hhe]r�F  (jdF  ]r�F  (h	he]r�F  (hh�e]r�F  (hhe]r�F  (jjF  ]r�F  (h	jlF  e]r�F  (hh�eeee]r�F  (hheeej�F  j�F  j�F  j�F  ]r�F  (jYF  ]r�F  (j[F  ]r�F  (j]F  ]r�F  (h	j_F  e]r�F  (hh�e]r�F  (hhe]r�F  (jdF  ]r�F  (h	he]r�F  (hh�e]r�F  (hhe]r�F  (jjF  ]r�F  (h	jlF  e]r�F  (hh�eeee]r�F  (hheeej�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  j�F  ]r�F  (jYF  ]r�F  (j[F  ]r�F  (j]F  ]r�F  (h	j_F  e]r G  (hh�e]rG  (hhe]rG  (jdF  ]rG  (h	he]rG  (hh�e]rG  (hhe]rG  (X	   Next-MoverG  ]rG  (h	h�e]r	G  (hh�eeee]r
G  (hheeej�F  j�F  j�F  j�F  j�F  j�F  ]rG  (jYF  ]rG  (j[F  ]rG  (j]F  ]rG  (h	j_F  e]rG  (hh�e]rG  (hhe]rG  (jdF  ]rG  (h	he]rG  (hh�e]rG  (hhe]rG  (jG  ]rG  (h	h�e]rG  (hh�eeee]rG  (hheee]rG  (jYF  ]rG  (j[F  ]rG  (j]F  ]rG  (h	j_F  e]rG  (hh�e]rG  (hhe]rG  (jdF  ]r G  (h	he]r!G  (hh�e]r"G  (hhe]r#G  (jG  ]r$G  (h	h�e]r%G  (hh�eeee]r&G  (hheeejG  jG  jG  jG  jG  jG  jG  jG  jG  jG  jG  jG  jG  jG  jG  ]r'G  (jYF  ]r(G  (j[F  ]r)G  (j]F  ]r*G  (h	j�  e]r+G  (hh�e]r,G  (hhe]r-G  (jdF  ]r.G  (h	he]r/G  (hh�e]r0G  (hhe]r1G  (jG  ]r2G  (h	h�e]r3G  (hh�eeee]r4G  (hheeej'G  j'G  ]r5G  (jYF  ]r6G  (j[F  ]r7G  (j]F  ]r8G  (h	j�  e]r9G  (hh�e]r:G  (hhe]r;G  (jdF  ]r<G  (h	he]r=G  (hh�e]r>G  (hhe]r?G  (jG  ]r@G  (h	h�e]rAG  (hh�eeee]rBG  (hheeej5G  ]rCG  (jYF  ]rDG  (j[F  ]rEG  (j]F  ]rFG  (h	j�  e]rGG  (hh�e]rHG  (hhe]rIG  (jdF  ]rJG  (h	he]rKG  (hh�e]rLG  (hhe]rMG  (jG  ]rNG  (h	h�e]rOG  (hh�eeee]rPG  (hheeejCG  jCG  jCG  jCG  ]rQG  (jYF  ]rRG  (j[F  ]rSG  (j]F  ]rTG  (h	j�  e]rUG  (hh�e]rVG  (hhe]rWG  (jdF  ]rXG  (h	he]rYG  (hh�e]rZG  (hhe]r[G  (jG  ]r\G  (h	h�e]r]G  (hh�eeee]r^G  (hheeejQG  jQG  jQG  jQG  jQG  jQG  jQG  jQG  jQG  jQG  ]r_G  (jYF  ]r`G  (j[F  ]raG  (j]F  ]rbG  (h	j�  e]rcG  (hh�e]rdG  (hhe]reG  (jdF  ]rfG  (h	he]rgG  (hh�e]rhG  (hhe]riG  (jG  ]rjG  (h	h�e]rkG  (hh�eeee]rlG  (hheeej_G  j_G  j_G  j_G  ]rmG  (jYF  ]rnG  (j[F  ]roG  (j]F  ]rpG  (h	j�  e]rqG  (hh�e]rrG  (hhe]rsG  (jdF  ]rtG  (h	he]ruG  (hh�e]rvG  (hhe]rwG  (jG  ]rxG  (h	h�e]ryG  (hh�eeee]rzG  (hheeejmG  jmG  ]r{G  (jYF  ]r|G  (j[F  ]r}G  (j]F  ]r~G  (h	j�  e]rG  (hh�e]r�G  (hhe]r�G  (jdF  ]r�G  (h	he]r�G  (hh�e]r�G  (hhe]r�G  (jG  ]r�G  (h	h�e]r�G  (hh�eeee]r�G  (hheeej{G  j{G  j{G  j{G  j{G  j{G  j{G  ]r�G  (jYF  ]r�G  (j[F  ]r�G  (j]F  ]r�G  (h	j�  e]r�G  (hh�e]r�G  (hhe]r�G  (jdF  ]r�G  (h	he]r�G  (hh�e]r�G  (hhe]r�G  (jG  ]r�G  (h	h�e]r�G  (hh�eeee]r�G  (hheee]r�G  (jYF  ]r�G  (j[F  ]r�G  (j]F  ]r�G  (h	j�  e]r�G  (hh�e]r�G  (hhe]r�G  (jdF  ]r�G  (h	he]r�G  (hh�e]r�G  (hhe]r�G  (jG  ]r�G  (h	h�e]r�G  (hh�eeee]r�G  (hheeej�G  ]r�G  (jYF  ]r�G  (j[F  ]r�G  (j]F  ]r�G  (h	j�  e]r�G  (hh�e]r�G  (hhe]r�G  (jdF  ]r�G  (h	he]r�G  (hh�e]r�G  (hhe]r�G  (jG  ]r�G  (h	h�e]r�G  (hh�eeee]r�G  (hheee]r�G  (jYF  ]r�G  (j[F  ]r�G  (j]F  ]r�G  (h	j�  e]r�G  (hh�e]r�G  (hhe]r�G  (jdF  ]r�G  (h	he]r�G  (hh�e]r�G  (hhe]r�G  (jG  ]r�G  (h	h�e]r�G  (hh�eeee]r�G  (hheeej�G  j�G  j�G  j�G  j�G  j�G  j�G  j�G  j�G  j�G  j�G  ]r�G  (jYF  ]r�G  (j[F  ]r�G  (j]F  ]r�G  (h	j�  e]r�G  (hh�e]r�G  (hhe]r�G  (jdF  ]r�G  (h	he]r�G  (hh�e]r�G  (hhe]r�G  (jG  ]r�G  (h	h�e]r�G  (hh�eeee]r�G  (hheeej�G  j�G  j�G  ]r�G  (jYF  ]r�G  (j[F  ]r�G  (j]F  ]r�G  (h	j�  e]r�G  (hh�e]r�G  (hhe]r�G  (jdF  ]r�G  (h	he]r�G  (hh�e]r�G  (hhe]r�G  (jG  ]r�G  (h	h�e]r�G  (hh�eeee]r�G  (hheeej�G  ]r�G  (jYF  ]r�G  (j[F  ]r�G  (j]F  ]r�G  (h	h�e]r�G  (hh�e]r�G  (hhe]r�G  (jdF  ]r�G  (h	he]r�G  (hh�e]r�G  (hhe]r�G  (jG  ]r�G  (h	h�e]r�G  (hh�eeee]r�G  (hheeej�G  ]r�G  (jYF  ]r�G  (j[F  ]r�G  (j]F  ]r�G  (h	h�e]r�G  (hh�e]r�G  (hhe]r�G  (jdF  ]r�G  (h	he]r�G  (hh�e]r�G  (hhe]r�G  (jG  ]r�G  (h	h�e]r�G  (hh�eeee]r�G  (hheee]r�G  (jYF  ]r�G  (j[F  ]r�G  (j]F  ]r�G  (h	h�e]r�G  (hh�e]r�G  (hhe]r�G  (jdF  ]r H  (h	he]rH  (hh�e]rH  (hhe]rH  (jG  ]rH  (h	h�e]rH  (hh�eeee]rH  (hheeej�G  ]rH  (jYF  ]rH  (j[F  ]r	H  (j]F  ]r
H  (h	h�e]rH  (hh�e]rH  (hhe]rH  (jdF  ]rH  (h	he]rH  (hh�e]rH  (hhe]rH  (jG  ]rH  (h	h�e]rH  (hh�eeee]rH  (hheeejH  ]rH  (jYF  ]rH  (j[F  ]rH  (j]F  ]rH  (h	h�e]rH  (hh�e]rH  (hhe]rH  (jdF  ]rH  (h	he]rH  (hh�e]rH  (hhe]rH  (jG  ]r H  (h	h�e]r!H  (hh�eeee]r"H  (hheeejH  ]r#H  (jYF  ]r$H  (j[F  ]r%H  (j]F  ]r&H  (h	h�e]r'H  (hh�e]r(H  (hhe]r)H  (jdF  ]r*H  (h	he]r+H  (hh�e]r,H  (hhe]r-H  (jG  ]r.H  (h	h�e]r/H  (hh�eeee]r0H  (hheeej#H  ]r1H  (jYF  ]r2H  (j[F  ]r3H  (j]F  ]r4H  (h	h�e]r5H  (hh�e]r6H  (hhe]r7H  (jdF  ]r8H  (h	he]r9H  (hh�e]r:H  (hhe]r;H  (jG  ]r<H  (h	h�e]r=H  (hh�eeee]r>H  (hheee]r?H  (jYF  ]r@H  (j[F  ]rAH  (j]F  ]rBH  (h	j�  e]rCH  (hh�e]rDH  (hhe]rEH  (jdF  ]rFH  (h	he]rGH  (hh�e]rHH  (hhe]rIH  (jG  ]rJH  (h	h�e]rKH  (hh�eeee]rLH  (hheeej?H  j?H  j?H  j?H  j?H  j?H  ]rMH  (jYF  ]rNH  (j[F  ]rOH  (j]F  ]rPH  (h	j�  e]rQH  (hh�e]rRH  (hhe]rSH  (jdF  ]rTH  (h	he]rUH  (hh�e]rVH  (hhe]rWH  (jG  ]rXH  (h	h�e]rYH  (hh�eeee]rZH  (hheeejMH  jMH  jMH  jMH  ]r[H  (jYF  ]r\H  (j[F  ]r]H  (j]F  ]r^H  (h	j�  e]r_H  (hh�e]r`H  (hhe]raH  (jdF  ]rbH  (h	he]rcH  (hh�e]rdH  (hhe]reH  (jG  ]rfH  (h	h�e]rgH  (hh�eeee]rhH  (hheee]riH  (jYF  ]rjH  (j[F  ]rkH  (j]F  ]rlH  (h	j�  e]rmH  (hh�e]rnH  (hhe]roH  (jdF  ]rpH  (h	he]rqH  (hh�e]rrH  (hhe]rsH  (jG  ]rtH  (h	h�e]ruH  (hh�eeee]rvH  (hheeejiH  jiH  jiH  jiH  jiH  jiH  jiH  jiH  jiH  ]rwH  (jYF  ]rxH  (j[F  ]ryH  (j]F  ]rzH  (h	j�  e]r{H  (hh�e]r|H  (hhe]r}H  (jdF  ]r~H  (h	he]rH  (hh�e]r�H  (hhe]r�H  (jG  ]r�H  (h	h�e]r�H  (hh�eeee]r�H  (hheee]r�H  (jYF  ]r�H  (j[F  ]r�H  (j]F  ]r�H  (h	j�  e]r�H  (hh�e]r�H  (hhe]r�H  (jdF  ]r�H  (h	he]r�H  (hh�e]r�H  (hhe]r�H  (jG  ]r�H  (h	h�e]r�H  (hh�eeee]r�H  (hheeej�H  j�H  ]r�H  (jYF  ]r�H  (j[F  ]r�H  (j]F  ]r�H  (h	j�  e]r�H  (hh�e]r�H  (hhe]r�H  (jdF  ]r�H  (h	he]r�H  (hh�e]r�H  (hhe]r�H  (jG  ]r�H  (h	h�e]r�H  (hh�eeee]r�H  (hheeej�H  ]r�H  (jYF  ]r�H  (j[F  ]r�H  (j]F  ]r�H  (h	j�  e]r�H  (hh�e]r�H  (hhe]r�H  (jdF  ]r�H  (h	he]r�H  (hh�e]r�H  (hhe]r�H  (jG  ]r�H  (h	h�e]r�H  (hh�eeee]r�H  (hheee]r�H  (jYF  ]r�H  (j[F  ]r�H  (j]F  ]r�H  (h	j�  e]r�H  (hh�e]r�H  (hhe]r�H  (jdF  ]r�H  (h	he]r�H  (hh�e]r�H  (hhe]r�H  (jG  ]r�H  (h	h�e]r�H  (hh�eeee]r�H  (hheeej�H  j�H  j�H  ]r�H  (jYF  ]r�H  (j[F  ]r�H  (j]F  ]r�H  (h	j�  e]r�H  (hh�e]r�H  (hhe]r�H  (jdF  ]r�H  (h	he]r�H  (hh�e]r�H  (hhe]r�H  (jG  ]r�H  (h	h�e]r�H  (hh�eeee]r�H  (hheee]r�H  (jYF  ]r�H  (j[F  ]r�H  (j]F  ]r�H  (h	j�  e]r�H  (hh�e]r�H  (hhe]r�H  (jdF  ]r�H  (h	he]r�H  (hh�e]r�H  (hhe]r�H  (jG  ]r�H  (h	h�e]r�H  (hh�eeee]r�H  (hheeej�H  ]r�H  (jYF  ]r�H  (j[F  ]r�H  (j]F  ]r�H  (h	j�  e]r�H  (hh�e]r�H  (hhe]r�H  (jdF  ]r�H  (h	he]r�H  (hh�e]r�H  (hhe]r�H  (jG  ]r�H  (h	h�e]r�H  (hh�eeee]r�H  (hheee]r�H  (jYF  ]r�H  (j[F  ]r�H  (j]F  ]r�H  (h	j�  e]r�H  (hh�e]r�H  (hhe]r�H  (jdF  ]r�H  (h	he]r�H  (hh�e]r�H  (hhe]r�H  (jG  ]r�H  (h	h�e]r�H  (hh�eeee]r�H  (hheeej�H  j�H  j�H  j�H  j�H  j�H  j�H  j�H  j�H  j�H  j�H  ]r�H  (jYF  ]r�H  (j[F  ]r�H  (j]F  ]r�H  (h	j�  e]r�H  (hh�e]r�H  (hhe]r�H  (jdF  ]r�H  (h	he]r�H  (hh�e]r�H  (hhe]r�H  (jG  ]r I  (h	h�e]rI  (hh�eeee]rI  (hheeej�H  j�H  j�H  ]rI  (jYF  ]rI  (j[F  ]rI  (j]F  ]rI  (h	j�  e]rI  (hh�e]rI  (hhe]r	I  (jdF  ]r
I  (h	he]rI  (hh�e]rI  (hhe]rI  (jG  ]rI  (h	h�e]rI  (hh�eeee]rI  (hheeejI  jI  ]rI  (jYF  ]rI  (j[F  ]rI  (j]F  ]rI  (h	j�  e]rI  (hh�e]rI  (hhe]rI  (jdF  ]rI  (h	he]rI  (hh�e]rI  (hhe]rI  (jG  ]rI  (h	h�e]rI  (hh�eeee]rI  (hheeejI  jI  jI  ]rI  (jYF  ]r I  (j[F  ]r!I  (j]F  ]r"I  (h	h�e]r#I  (hh�e]r$I  (hhe]r%I  (jdF  ]r&I  (h	he]r'I  (hh�e]r(I  (hhe]r)I  (jG  ]r*I  (h	h�e]r+I  (hh�eeee]r,I  (hheee]r-I  (jYF  ]r.I  (j[F  ]r/I  (j]F  ]r0I  (h	h�e]r1I  (hh�e]r2I  (hhe]r3I  (jdF  ]r4I  (h	he]r5I  (hh�e]r6I  (hhe]r7I  (jG  ]r8I  (h	h�e]r9I  (hh�eeee]r:I  (hheeej-I  j-I  j-I  j-I  j-I  j-I  j-I  j-I  j-I  j-I  j-I  j-I  j-I  j-I  j-I  j-I  ]r;I  (jYF  ]r<I  (j[F  ]r=I  (j]F  ]r>I  (h	h�e]r?I  (hh�e]r@I  (hhe]rAI  (jdF  ]rBI  (h	he]rCI  (hh�e]rDI  (hhe]rEI  (jG  ]rFI  (h	h�e]rGI  (hh�eeee]rHI  (hheeej;I  j;I  j;I  j;I  ]rII  (jYF  ]rJI  (j[F  ]rKI  (j]F  ]rLI  (h	h�e]rMI  (hh�e]rNI  (hhe]rOI  (jdF  ]rPI  (h	he]rQI  (hh�e]rRI  (hhe]rSI  (jG  ]rTI  (h	h�e]rUI  (hh�eeee]rVI  (hheeejII  ]rWI  (jYF  ]rXI  (j[F  ]rYI  (j]F  ]rZI  (h	h�e]r[I  (hh�e]r\I  (hhe]r]I  (jdF  ]r^I  (h	he]r_I  (hh�e]r`I  (hhe]raI  (jG  ]rbI  (h	h�e]rcI  (hh�eeee]rdI  (hheee]reI  (jYF  ]rfI  (j[F  ]rgI  (j]F  ]rhI  (h	h�e]riI  (hh�e]rjI  (hhe]rkI  (jdF  ]rlI  (h	he]rmI  (hh�e]rnI  (hhe]roI  (jG  ]rpI  (h	h�e]rqI  (hh�eeee]rrI  (hheeejeI  ]rsI  (jYF  ]rtI  (j[F  ]ruI  (j]F  ]rvI  (h	h�e]rwI  (hh�e]rxI  (hhe]ryI  (jdF  ]rzI  (h	he]r{I  (hh�e]r|I  (hhe]r}I  (jG  ]r~I  (h	h�e]rI  (hh�eeee]r�I  (hheeejsI  jsI  jsI  jsI  jsI  ]r�I  (jYF  ]r�I  (j[F  ]r�I  (j]F  ]r�I  (h	h�e]r�I  (hh�e]r�I  (hhe]r�I  (jdF  ]r�I  (h	he]r�I  (hh�e]r�I  (hhe]r�I  (jG  ]r�I  (h	h�e]r�I  (hh�eeee]r�I  (hheeej�I  ]r�I  (jYF  ]r�I  (j[F  ]r�I  (j]F  ]r�I  (h	h�e]r�I  (hh�e]r�I  (hhe]r�I  (jdF  ]r�I  (h	he]r�I  (hh�e]r�I  (hhe]r�I  (jG  ]r�I  (h	h�e]r�I  (hh�eeee]r�I  (hheeej�I  ]r�I  (jYF  ]r�I  (j[F  ]r�I  (j]F  ]r�I  (h	h�e]r�I  (hh�e]r�I  (hhe]r�I  (jdF  ]r�I  (h	he]r�I  (hh�e]r�I  (hhe]r�I  (jG  ]r�I  (h	h�e]r�I  (hh�eeee]r�I  (hheee]r�I  (jYF  ]r�I  (j[F  ]r�I  (j]F  ]r�I  (h	h�e]r�I  (hh�e]r�I  (hhe]r�I  (jdF  ]r�I  (h	he]r�I  (hh�e]r�I  (hhe]r�I  (jG  ]r�I  (h	h�e]r�I  (hh�eeee]r�I  (hheeej�I  j�I  j�I  j�I  ]r�I  (jYF  ]r�I  (j[F  ]r�I  (j]F  ]r�I  (h	h�e]r�I  (hh�e]r�I  (hhe]r�I  (jdF  ]r�I  (h	he]r�I  (hh�e]r�I  (hhe]r�I  (jG  ]r�I  (h	h�e]r�I  (hh�eeee]r�I  (hheeej�I  j�I  j�I  j�I  ]r�I  (jYF  ]r�I  (j[F  ]r�I  (j]F  ]r�I  (h	h�e]r�I  (hh�e]r�I  (hhe]r�I  (jdF  ]r�I  (h	he]r�I  (hh�e]r�I  (hhe]r�I  (jG  ]r�I  (h	h�e]r�I  (hh�eeee]r�I  (hheeej�I  j�I  j�I  j�I  j�I  j�I  j�I  ]r�I  (jYF  ]r�I  (j[F  ]r�I  (j]F  ]r�I  (h	h�e]r�I  (hh�e]r�I  (hhe]r�I  (jdF  ]r�I  (h	he]r�I  (hh�e]r�I  (hhe]r�I  (jG  ]r�I  (h	h�e]r�I  (hh�eeee]r�I  (hheeej�I  j�I  j�I  j�I  ]r�I  (jYF  ]r�I  (j[F  ]r�I  (j]F  ]r�I  (h	h�e]r�I  (hh�e]r�I  (hhe]r�I  (jdF  ]r�I  (h	he]r�I  (hh�e]r�I  (hhe]r�I  (jG  ]r�I  (h	h�e]r�I  (hh�eeee]r�I  (hheeej�I  ]r�I  (jYF  ]r�I  (j[F  ]r�I  (j]F  ]r�I  (h	h�e]r�I  (hh�e]r�I  (hhe]r�I  (jdF  ]r�I  (h	he]r�I  (hh�e]r�I  (hhe]r�I  (jG  ]r�I  (h	h�e]r�I  (hh�eeee]r�I  (hheee]r�I  (jYF  ]r J  (j[F  ]rJ  (j]F  ]rJ  (h	h�e]rJ  (hh�e]rJ  (hhe]rJ  (jdF  ]rJ  (h	he]rJ  (hh�e]rJ  (hhe]r	J  (jG  ]r
J  (h	h�e]rJ  (hh�eeee]rJ  (hheeej�I  j�I  j�I  j�I  j�I  j�I  j�I  ]rJ  (jYF  ]rJ  (j[F  ]rJ  (j]F  ]rJ  (h	h�e]rJ  (hh�e]rJ  (hhe]rJ  (jdF  ]rJ  (h	he]rJ  (hh�e]rJ  (hhe]rJ  (jG  ]rJ  (h	h�e]rJ  (hh�eeee]rJ  (hheeejJ  jJ  jJ  jJ  ]rJ  (jYF  ]rJ  (j[F  ]rJ  (j]F  ]rJ  (h	h�e]rJ  (hh�e]r J  (hhe]r!J  (jdF  ]r"J  (h	he]r#J  (hh�e]r$J  (hhe]r%J  (jG  ]r&J  (h	h�e]r'J  (hh�eeee]r(J  (hheee]r)J  (jYF  ]r*J  (j[F  ]r+J  (j]F  ]r,J  (h	h�e]r-J  (hh�e]r.J  (hhe]r/J  (jdF  ]r0J  (h	he]r1J  (hh�e]r2J  (hhe]r3J  (jG  ]r4J  (h	h�e]r5J  (hh�eeee]r6J  (hheeej)J  ]r7J  (jYF  ]r8J  (j[F  ]r9J  (j]F  ]r:J  (h	h�e]r;J  (hh�e]r<J  (hhe]r=J  (jdF  ]r>J  (h	he]r?J  (hh�e]r@J  (hhe]rAJ  (jG  ]rBJ  (h	h�e]rCJ  (hh�eeee]rDJ  (hheeej7J  j7J  ]rEJ  (jYF  ]rFJ  (j[F  ]rGJ  (j]F  ]rHJ  (h	h�e]rIJ  (hh�e]rJJ  (hhe]rKJ  (jdF  ]rLJ  (h	he]rMJ  (hh�e]rNJ  (hhe]rOJ  (jG  ]rPJ  (h	h�e]rQJ  (hh�eeee]rRJ  (hheee]rSJ  (jYF  ]rTJ  (j[F  ]rUJ  (j]F  ]rVJ  (h	h�e]rWJ  (hh�e]rXJ  (hhe]rYJ  (jdF  ]rZJ  (h	he]r[J  (hh�e]r\J  (hhe]r]J  (jG  ]r^J  (h	h�e]r_J  (hh�eeee]r`J  (hheeejSJ  ]raJ  (jYF  ]rbJ  (j[F  ]rcJ  (j]F  ]rdJ  (h	h�e]reJ  (hh�e]rfJ  (hhe]rgJ  (jdF  ]rhJ  (h	he]riJ  (hh�e]rjJ  (hhe]rkJ  (jG  ]rlJ  (h	h�e]rmJ  (hh�eeee]rnJ  (hheeejaJ  ]roJ  (jYF  ]rpJ  (j[F  ]rqJ  (j]F  ]rrJ  (h	h�e]rsJ  (hh�e]rtJ  (hhe]ruJ  (jdF  ]rvJ  (h	he]rwJ  (hh�e]rxJ  (hhe]ryJ  (jG  ]rzJ  (h	h�e]r{J  (hh�eeee]r|J  (hheeejoJ  joJ  joJ  joJ  joJ  ]r}J  (jYF  ]r~J  (j[F  ]rJ  (j]F  ]r�J  (h	h�e]r�J  (hh�e]r�J  (hhe]r�J  (jdF  ]r�J  (h	he]r�J  (hh�e]r�J  (hhe]r�J  (jG  ]r�J  (h	h�e]r�J  (hh�eeee]r�J  (hheeej}J  ]r�J  (jYF  ]r�J  (j[F  ]r�J  (j]F  ]r�J  (h	h�e]r�J  (hh�e]r�J  (hhe]r�J  (jdF  ]r�J  (h	he]r�J  (hh�e]r�J  (hhe]r�J  (jG  ]r�J  (h	h�e]r�J  (hh�eeee]r�J  (hheeej�J  ]r�J  (jYF  ]r�J  (j[F  ]r�J  (j]F  ]r�J  (h	h�e]r�J  (hh�e]r�J  (hhe]r�J  (jdF  ]r�J  (h	he]r�J  (hh�e]r�J  (hhe]r�J  (jG  ]r�J  (h	h�e]r�J  (hh�eeee]r�J  (hheeej�J  j�J  j�J  j�J  ]r�J  (jYF  ]r�J  (j[F  ]r�J  (j]F  ]r�J  (h	h�e]r�J  (hh�e]r�J  (hhe]r�J  (jdF  ]r�J  (h	he]r�J  (hh�e]r�J  (hhe]r�J  (jG  ]r�J  (h	h�e]r�J  (hh�eeee]r�J  (hheeej�J  j�J  j�J  j�J  j�J  j�J  j�J  j�J  j�J  j�J  j�J  j�J  ]r�J  (jYF  ]r�J  (j[F  ]r�J  (j]F  ]r�J  (h	h�e]r�J  (hh�e]r�J  (hhe]r�J  (jdF  ]r�J  (h	he]r�J  (hh�e]r�J  (hhe]r�J  (jG  ]r�J  (h	h�e]r�J  (hh�eeee]r�J  (hheeej�J  j�J  j�J  j�J  j�J  ]r�J  (jYF  ]r�J  (j[F  ]r�J  (j]F  ]r�J  (h	h�e]r�J  (hh�e]r�J  (hhe]r�J  (jdF  ]r�J  (h	he]r�J  (hh�e]r�J  (hhe]r�J  (jG  ]r�J  (h	h�e]r�J  (hh�eeee]r�J  (hheeej�J  ]r�J  (jYF  ]r�J  (j[F  ]r�J  (j]F  ]r�J  (h	h�e]r�J  (hh�e]r�J  (hhe]r�J  (jdF  ]r�J  (h	he]r�J  (hh�e]r�J  (hhe]r�J  (jG  ]r�J  (h	h�e]r�J  (hh�eeee]r�J  (hheeej�J  j�J  ]r�J  (jYF  ]r�J  (j[F  ]r�J  (j]F  ]r�J  (h	h�e]r�J  (hh�e]r�J  (hhe]r�J  (jdF  ]r�J  (h	he]r�J  (hh�e]r�J  (hhe]r�J  (jG  ]r�J  (h	h�e]r�J  (hh�eeee]r�J  (hheeej�J  j�J  j�J  j�J  j�J  j�J  ]r�J  (jYF  ]r�J  (j[F  ]r�J  (j]F  ]r�J  (h	h�e]r�J  (hh�e]r�J  (hhe]r�J  (jdF  ]r�J  (h	he]r�J  (hh�e]r�J  (hhe]r�J  (jG  ]r�J  (h	h�e]r�J  (hh�eeee]r�J  (hheee]r�J  (jYF  ]r�J  (j[F  ]r�J  (j]F  ]r�J  (h	h�e]r�J  (hh�e]r K  (hhe]rK  (jdF  ]rK  (h	he]rK  (hh�e]rK  (hhe]rK  (jG  ]rK  (h	h�e]rK  (hh�eeee]rK  (hheeej�J  j�J  ]r	K  (jYF  ]r
K  (j[F  ]rK  (j]F  ]rK  (h	h�e]rK  (hh�e]rK  (hhe]rK  (jdF  ]rK  (h	he]rK  (hh�e]rK  (hhe]rK  (jG  ]rK  (h	h�e]rK  (hh�eeee]rK  (hheeej	K  j	K  j	K  j	K  j	K  j	K  j	K  ]rK  (jYF  ]rK  (j[F  ]rK  (j]F  ]rK  (h	h�e]rK  (hh�e]rK  (hhe]rK  (jdF  ]rK  (h	he]rK  (hh�e]r K  (hhe]r!K  (jG  ]r"K  (h	h�e]r#K  (hh�eeee]r$K  (hheee]r%K  (jYF  ]r&K  (j[F  ]r'K  (j]F  ]r(K  (h	h�e]r)K  (hh�e]r*K  (hhe]r+K  (jdF  ]r,K  (h	he]r-K  (hh�e]r.K  (hhe]r/K  (jG  ]r0K  (h	h�e]r1K  (hh�eeee]r2K  (hheeej%K  j%K  j%K  j%K  j%K  j%K  j%K  j%K  j%K  j%K  ]r3K  (jYF  ]r4K  (j[F  ]r5K  (j]F  ]r6K  (h	h�e]r7K  (hh�e]r8K  (hhe]r9K  (jdF  ]r:K  (h	he]r;K  (hh�e]r<K  (hhe]r=K  (jG  ]r>K  (h	h�e]r?K  (hh�eeee]r@K  (hheeej3K  ]rAK  (jYF  ]rBK  (j[F  ]rCK  (j]F  ]rDK  (h	h�e]rEK  (hh�e]rFK  (hhe]rGK  (jdF  ]rHK  (h	he]rIK  (hh�e]rJK  (hhe]rKK  (jG  ]rLK  (h	h�e]rMK  (hh�eeee]rNK  (hheeejAK  ]rOK  (jYF  ]rPK  (j[F  ]rQK  (j]F  ]rRK  (h	h�e]rSK  (hh�e]rTK  (hhe]rUK  (jdF  ]rVK  (h	he]rWK  (hh�e]rXK  (hhe]rYK  (jG  ]rZK  (h	h�e]r[K  (hh�eeee]r\K  (hheeejOK  ]r]K  (jYF  ]r^K  (j[F  ]r_K  (j]F  ]r`K  (h	h�e]raK  (hh�e]rbK  (hhe]rcK  (jdF  ]rdK  (h	he]reK  (hh�e]rfK  (hhe]rgK  (jG  ]rhK  (h	h�e]riK  (hh�eeee]rjK  (hheee]rkK  (jYF  ]rlK  (j[F  ]rmK  (j]F  ]rnK  (h	j�  e]roK  (hh�e]rpK  (hhe]rqK  (jdF  ]rrK  (h	he]rsK  (hh�e]rtK  (hhe]ruK  (jG  ]rvK  (h	h�e]rwK  (hh�eeee]rxK  (hheee]ryK  (jYF  ]rzK  (j[F  ]r{K  (j]F  ]r|K  (h	j�  e]r}K  (hh�e]r~K  (hhe]rK  (jdF  ]r�K  (h	he]r�K  (hh�e]r�K  (hhe]r�K  (jG  ]r�K  (h	h�e]r�K  (hh�eeee]r�K  (hheeejyK  ]r�K  (jYF  ]r�K  (j[F  ]r�K  (j]F  ]r�K  (h	j�  e]r�K  (hh�e]r�K  (hhe]r�K  (jdF  ]r�K  (h	he]r�K  (hh�e]r�K  (hhe]r�K  (jG  ]r�K  (h	h�e]r�K  (hh�eeee]r�K  (hheeej�K  j�K  j�K  j�K  j�K  j�K  ]r�K  (jYF  ]r�K  (j[F  ]r�K  (j]F  ]r�K  (h	j�  e]r�K  (hh�e]r�K  (hhe]r�K  (jdF  ]r�K  (h	he]r�K  (hh�e]r�K  (hhe]r�K  (jG  ]r�K  (h	h�e]r�K  (hh�eeee]r�K  (hheeej�K  j�K  ]r�K  (jYF  ]r�K  (j[F  ]r�K  (j]F  ]r�K  (h	j�  e]r�K  (hh�e]r�K  (hhe]r�K  (jdF  ]r�K  (h	he]r�K  (hh�e]r�K  (hhe]r�K  (jG  ]r�K  (h	h�e]r�K  (hh�eeee]r�K  (hheee]r�K  (jYF  ]r�K  (j[F  ]r�K  (j]F  ]r�K  (h	j�  e]r�K  (hh�e]r�K  (hhe]r�K  (jdF  ]r�K  (h	he]r�K  (hh�e]r�K  (hhe]r�K  (jG  ]r�K  (h	h�e]r�K  (hh�eeee]r�K  (hheeej�K  j�K  j�K  j�K  j�K  j�K  j�K  j�K  ]r�K  (jYF  ]r�K  (j[F  ]r�K  (j]F  ]r�K  (h	j�  e]r�K  (hh�e]r�K  (hhe]r�K  (jdF  ]r�K  (h	he]r�K  (hh�e]r�K  (hhe]r�K  (jG  ]r�K  (h	h�e]r�K  (hh�eeee]r�K  (hheee]r�K  (jYF  ]r�K  (j[F  ]r�K  (j]F  ]r�K  (h	j�  e]r�K  (hh�e]r�K  (hhe]r�K  (jdF  ]r�K  (h	he]r�K  (hh�e]r�K  (hhe]r�K  (jG  ]r�K  (h	h�e]r�K  (hh�eeee]r�K  (hheeej�K  j�K  j�K  j�K  j�K  ]r�K  (jYF  ]r�K  (j[F  ]r�K  (j]F  ]r�K  (h	j�  e]r�K  (hh�e]r�K  (hhe]r�K  (jdF  ]r�K  (h	he]r�K  (hh�e]r�K  (hhe]r�K  (X	   Next-Mover�K  ]r�K  (h	h�e]r�K  (hh�eeee]r�K  (hheeej�K  j�K  ]r�K  (jYF  ]r�K  (j[F  ]r�K  (j]F  ]r�K  (h	j�  e]r�K  (hh�e]r�K  (hhe]r�K  (jdF  ]r�K  (h	he]r�K  (hh�e]r�K  (hhe]r�K  (j�K  ]r�K  (h	h�e]r�K  (hh�eeee]r�K  (hheee]r�K  (jYF  ]r�K  (j[F  ]r�K  (j]F  ]r�K  (h	j�  e]r�K  (hh�e]r�K  (hhe]r�K  (jdF  ]r�K  (h	he]r L  (hh�e]rL  (hhe]rL  (j�K  ]rL  (h	h�e]rL  (hh�eeee]rL  (hheee]rL  (jYF  ]rL  (j[F  ]rL  (j]F  ]r	L  (h	j�  e]r
L  (hh�e]rL  (hhe]rL  (jdF  ]rL  (h	he]rL  (hh�e]rL  (hhe]rL  (j�K  ]rL  (h	h�e]rL  (hh�eeee]rL  (hheeejL  jL  jL  jL  jL  jL  jL  jL  jL  jL  jL  jL  jL  jL  jL  jL  jL  jL  jL  jL  jL  ]rL  (jYF  ]rL  (j[F  ]rL  (j]F  ]rL  (h	j�  e]rL  (hh�e]rL  (hhe]rL  (jdF  ]rL  (h	he]rL  (hh�e]rL  (hhe]rL  (j�K  ]rL  (h	h�e]r L  (hh�eeee]r!L  (hheeejL  jL  jL  jL  jL  jL  ]r"L  (jYF  ]r#L  (j[F  ]r$L  (j]F  ]r%L  (h	j�  e]r&L  (hh�e]r'L  (hhe]r(L  (jdF  ]r)L  (h	he]r*L  (hh�e]r+L  (hhe]r,L  (j�K  ]r-L  (h	h�e]r.L  (hh�eeee]r/L  (hheee]r0L  (jYF  ]r1L  (j[F  ]r2L  (j]F  ]r3L  (h	j�  e]r4L  (hh�e]r5L  (hhe]r6L  (jdF  ]r7L  (h	he]r8L  (hh�e]r9L  (hhe]r:L  (j�K  ]r;L  (h	h�e]r<L  (hh�eeee]r=L  (hheee]r>L  (jYF  ]r?L  (j[F  ]r@L  (j]F  ]rAL  (h	j�  e]rBL  (hh�e]rCL  (hhe]rDL  (jdF  ]rEL  (h	he]rFL  (hh�e]rGL  (hhe]rHL  (j�K  ]rIL  (h	h�e]rJL  (hh�eeee]rKL  (hheeej>L  ]rLL  (jYF  ]rML  (j[F  ]rNL  (j]F  ]rOL  (h	j�  e]rPL  (hh�e]rQL  (hhe]rRL  (jdF  ]rSL  (h	he]rTL  (hh�e]rUL  (hhe]rVL  (j�K  ]rWL  (h	h�e]rXL  (hh�eeee]rYL  (hheeejLL  jLL  jLL  jLL  jLL  ]rZL  (jYF  ]r[L  (j[F  ]r\L  (j]F  ]r]L  (h	j�  e]r^L  (hh�e]r_L  (hhe]r`L  (jdF  ]raL  (h	he]rbL  (hh�e]rcL  (hhe]rdL  (j�K  ]reL  (h	h�e]rfL  (hh�eeee]rgL  (hheeejZL  jZL  jZL  ]rhL  (jYF  ]riL  (j[F  ]rjL  (j]F  ]rkL  (h	j�  e]rlL  (hh�e]rmL  (hhe]rnL  (jdF  ]roL  (h	he]rpL  (hh�e]rqL  (hhe]rrL  (j�K  ]rsL  (h	h�e]rtL  (hh�eeee]ruL  (hheee]rvL  (jYF  ]rwL  (j[F  ]rxL  (j]F  ]ryL  (h	j�  e]rzL  (hh�e]r{L  (hhe]r|L  (jdF  ]r}L  (h	he]r~L  (hh�e]rL  (hhe]r�L  (j�K  ]r�L  (h	h�e]r�L  (hh�eeee]r�L  (hheeejvL  jvL  jvL  jvL  ]r�L  (jYF  ]r�L  (j[F  ]r�L  (j]F  ]r�L  (h	j�  e]r�L  (hh�e]r�L  (hhe]r�L  (jdF  ]r�L  (h	he]r�L  (hh�e]r�L  (hhe]r�L  (j�K  ]r�L  (h	h�e]r�L  (hh�eeee]r�L  (hheee]r�L  (jYF  ]r�L  (j[F  ]r�L  (j]F  ]r�L  (h	j�  e]r�L  (hh�e]r�L  (hhe]r�L  (jdF  ]r�L  (h	he]r�L  (hh�e]r�L  (hhe]r�L  (j�K  ]r�L  (h	h�e]r�L  (hh�eeee]r�L  (hheeej�L  j�L  j�L  j�L  j�L  ]r�L  (jYF  ]r�L  (j[F  ]r�L  (j]F  ]r�L  (h	j�  e]r�L  (hh�e]r�L  (hhe]r�L  (jdF  ]r�L  (h	he]r�L  (hh�e]r�L  (hhe]r�L  (j�K  ]r�L  (h	h�e]r�L  (hh�eeee]r�L  (hheeej�L  j�L  j�L  ]r�L  (jYF  ]r�L  (j[F  ]r�L  (j]F  ]r�L  (h	j�  e]r�L  (hh�e]r�L  (hhe]r�L  (jdF  ]r�L  (h	he]r�L  (hh�e]r�L  (hhe]r�L  (j�K  ]r�L  (h	h�e]r�L  (hh�eeee]r�L  (hheeej�L  ]r�L  (jYF  ]r�L  (j[F  ]r�L  (j]F  ]r�L  (h	j�  e]r�L  (hh�e]r�L  (hhe]r�L  (jdF  ]r�L  (h	he]r�L  (hh�e]r�L  (hhe]r�L  (j�K  ]r�L  (h	h�e]r�L  (hh�eeee]r�L  (hheeej�L  ]r�L  (jYF  ]r�L  (j[F  ]r�L  (j]F  ]r�L  (h	j�  e]r�L  (hh�e]r�L  (hhe]r�L  (jdF  ]r�L  (h	he]r�L  (hh�e]r�L  (hhe]r�L  (j�K  ]r�L  (h	h�e]r�L  (hh�eeee]r�L  (hheeej�L  j�L  ]r�L  (jYF  ]r�L  (j[F  ]r�L  (j]F  ]r�L  (h	j�  e]r�L  (hh�e]r�L  (hhe]r�L  (jdF  ]r�L  (h	he]r�L  (hh�e]r�L  (hhe]r�L  (j�K  ]r�L  (h	h�e]r�L  (hh�eeee]r�L  (hheeej�L  j�L  j�L  ]r�L  (jYF  ]r�L  (j[F  ]r�L  (j]F  ]r�L  (h	j�  e]r�L  (hh�e]r�L  (hhe]r�L  (jdF  ]r�L  (h	he]r�L  (hh�e]r�L  (hhe]r�L  (j�K  ]r�L  (h	h�e]r�L  (hh�eeee]r�L  (hheeej�L  j�L  j�L  j�L  ]r�L  (jYF  ]r�L  (j[F  ]r�L  (j]F  ]r�L  (h	j�  e]r�L  (hh�e]r�L  (hhe]r�L  (jdF  ]r�L  (h	he]r�L  (hh�e]r�L  (hhe]r�L  (j�K  ]r�L  (h	h�e]r M  (hh�eeee]rM  (hheeej�L  ]rM  (jYF  ]rM  (j[F  ]rM  (j]F  ]rM  (h	j�  e]rM  (hh�e]rM  (hhe]rM  (jdF  ]r	M  (h	he]r
M  (hh�e]rM  (hhe]rM  (j�K  ]rM  (h	h�e]rM  (hh�eeee]rM  (hheeejM  jM  jM  jM  ]rM  (jYF  ]rM  (j[F  ]rM  (j]F  ]rM  (h	j�  e]rM  (hh�e]rM  (hhe]rM  (jdF  ]rM  (h	he]rM  (hh�e]rM  (hhe]rM  (j�K  ]rM  (h	h�e]rM  (hh�eeee]rM  (hheeejM  jM  ]rM  (jYF  ]rM  (j[F  ]r M  (j]F  ]r!M  (h	j�  e]r"M  (hh�e]r#M  (hhe]r$M  (jdF  ]r%M  (h	he]r&M  (hh�e]r'M  (hhe]r(M  (j�K  ]r)M  (h	h�e]r*M  (hh�eeee]r+M  (hheeejM  jM  ]r,M  (jYF  ]r-M  (j[F  ]r.M  (j]F  ]r/M  (h	j�  e]r0M  (hh�e]r1M  (hhe]r2M  (jdF  ]r3M  (h	he]r4M  (hh�e]r5M  (hhe]r6M  (j�K  ]r7M  (h	h�e]r8M  (hh�eeee]r9M  (hheeej,M  ]r:M  (jYF  ]r;M  (j[F  ]r<M  (j]F  ]r=M  (h	j�  e]r>M  (hh�e]r?M  (hhe]r@M  (jdF  ]rAM  (h	he]rBM  (hh�e]rCM  (hhe]rDM  (j�K  ]rEM  (h	h�e]rFM  (hh�eeee]rGM  (hheeej:M  j:M  j:M  ]rHM  (jYF  ]rIM  (j[F  ]rJM  (j]F  ]rKM  (h	j�  e]rLM  (hh�e]rMM  (hhe]rNM  (jdF  ]rOM  (h	he]rPM  (hh�e]rQM  (hhe]rRM  (j�K  ]rSM  (h	h�e]rTM  (hh�eeee]rUM  (hheeejHM  jHM  jHM  jHM  jHM  ]rVM  (jYF  ]rWM  (j[F  ]rXM  (j]F  ]rYM  (h	j�  e]rZM  (hh�e]r[M  (hhe]r\M  (jdF  ]r]M  (h	he]r^M  (hh�e]r_M  (hhe]r`M  (j�K  ]raM  (h	h�e]rbM  (hh�eeee]rcM  (hheee]rdM  (jYF  ]reM  (j[F  ]rfM  (j]F  ]rgM  (h	j�  e]rhM  (hh�e]riM  (hhe]rjM  (jdF  ]rkM  (h	he]rlM  (hh�e]rmM  (hhe]rnM  (j�K  ]roM  (h	h�e]rpM  (hh�eeee]rqM  (hheeejdM  jdM  jdM  jdM  ]rrM  (jYF  ]rsM  (j[F  ]rtM  (j]F  ]ruM  (h	j�  e]rvM  (hh�e]rwM  (hhe]rxM  (jdF  ]ryM  (h	he]rzM  (hh�e]r{M  (hhe]r|M  (j�K  ]r}M  (h	h�e]r~M  (hh�eeee]rM  (hheeejrM  jrM  ]r�M  (jYF  ]r�M  (j[F  ]r�M  (j]F  ]r�M  (h	j�  e]r�M  (hh�e]r�M  (hhe]r�M  (jdF  ]r�M  (h	he]r�M  (hh�e]r�M  (hhe]r�M  (j�K  ]r�M  (h	h�e]r�M  (hh�eeee]r�M  (hheeej�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  ]r�M  (jYF  ]r�M  (j[F  ]r�M  (j]F  ]r�M  (h	j�  e]r�M  (hh�e]r�M  (hhe]r�M  (jdF  ]r�M  (h	he]r�M  (hh�e]r�M  (hhe]r�M  (j�K  ]r�M  (h	h�e]r�M  (hh�eeee]r�M  (hheeej�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  ]r�M  (jYF  ]r�M  (j[F  ]r�M  (j]F  ]r�M  (h	j�  e]r�M  (hh�e]r�M  (hhe]r�M  (jdF  ]r�M  (h	he]r�M  (hh�e]r�M  (hhe]r�M  (j�K  ]r�M  (h	h�e]r�M  (hh�eeee]r�M  (hheeej�M  j�M  j�M  ]r�M  (jYF  ]r�M  (j[F  ]r�M  (j]F  ]r�M  (h	j�  e]r�M  (hh�e]r�M  (hhe]r�M  (jdF  ]r�M  (h	he]r�M  (hh�e]r�M  (hhe]r�M  (j�K  ]r�M  (h	h�e]r�M  (hh�eeee]r�M  (hheee]r�M  (jYF  ]r�M  (j[F  ]r�M  (j]F  ]r�M  (h	j�  e]r�M  (hh�e]r�M  (hhe]r�M  (jdF  ]r�M  (h	he]r�M  (hh�e]r�M  (hhe]r�M  (j�K  ]r�M  (h	h�e]r�M  (hh�eeee]r�M  (hheee]r�M  (jYF  ]r�M  (j[F  ]r�M  (j]F  ]r�M  (h	j�  e]r�M  (hh�e]r�M  (hhe]r�M  (jdF  ]r�M  (h	he]r�M  (hh�e]r�M  (hhe]r�M  (j�K  ]r�M  (h	h�e]r�M  (hh�eeee]r�M  (hheeej�M  j�M  j�M  j�M  j�M  ]r�M  (jYF  ]r�M  (j[F  ]r�M  (j]F  ]r�M  (h	j�  e]r�M  (hh�e]r�M  (hhe]r�M  (jdF  ]r�M  (h	he]r�M  (hh�e]r�M  (hhe]r�M  (j�K  ]r�M  (h	h�e]r�M  (hh�eeee]r�M  (hheeej�M  ]r�M  (jYF  ]r�M  (j[F  ]r�M  (j]F  ]r�M  (h	j�  e]r�M  (hh�e]r�M  (hhe]r�M  (jdF  ]r�M  (h	he]r�M  (hh�e]r�M  (hhe]r�M  (j�K  ]r�M  (h	h�e]r�M  (hh�eeee]r�M  (hheee]r�M  (jYF  ]r�M  (j[F  ]r�M  (j]F  ]r�M  (h	j�  e]r�M  (hh�e]r�M  (hhe]r�M  (jdF  ]r�M  (h	he]r�M  (hh�e]r�M  (hhe]r�M  (j�K  ]r�M  (h	h�e]r�M  (hh�eeee]r�M  (hheee]r�M  (jYF  ]r�M  (j[F  ]r N  (j]F  ]rN  (h	j�  e]rN  (hh�e]rN  (hhe]rN  (jdF  ]rN  (h	he]rN  (hh�e]rN  (hhe]rN  (j�K  ]r	N  (h	h�e]r
N  (hh�eeee]rN  (hheeej�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  j�M  ]rN  (jYF  ]rN  (j[F  ]rN  (j]F  ]rN  (h	h�e]rN  (hh�e]rN  (hhe]rN  (jdF  ]rN  (h	he]rN  (hh�e]rN  (hhe]rN  (j�K  ]rN  (h	h�e]rN  (hh�eeee]rN  (hheeejN  ]rN  (jYF  ]rN  (j[F  ]rN  (j]F  ]rN  (h	h�e]rN  (hh�e]rN  (hhe]r N  (jdF  ]r!N  (h	he]r"N  (hh�e]r#N  (hhe]r$N  (j�K  ]r%N  (h	h�e]r&N  (hh�eeee]r'N  (hheeejN  ]r(N  (jYF  ]r)N  (j[F  ]r*N  (j]F  ]r+N  (h	h�e]r,N  (hh�e]r-N  (hhe]r.N  (jdF  ]r/N  (h	he]r0N  (hh�e]r1N  (hhe]r2N  (j�K  ]r3N  (h	h�e]r4N  (hh�eeee]r5N  (hheeej(N  j(N  j(N  ]r6N  (jYF  ]r7N  (j[F  ]r8N  (j]F  ]r9N  (h	h�e]r:N  (hh�e]r;N  (hhe]r<N  (jdF  ]r=N  (h	he]r>N  (hh�e]r?N  (hhe]r@N  (j�K  ]rAN  (h	h�e]rBN  (hh�eeee]rCN  (hheeej6N  j6N  ]rDN  (jYF  ]rEN  (j[F  ]rFN  (j]F  ]rGN  (h	h�e]rHN  (hh�e]rIN  (hhe]rJN  (jdF  ]rKN  (h	he]rLN  (hh�e]rMN  (hhe]rNN  (j�K  ]rON  (h	h�e]rPN  (hh�eeee]rQN  (hheeejDN  ]rRN  (jYF  ]rSN  (j[F  ]rTN  (j]F  ]rUN  (h	h�e]rVN  (hh�e]rWN  (hhe]rXN  (jdF  ]rYN  (h	he]rZN  (hh�e]r[N  (hhe]r\N  (j�K  ]r]N  (h	h�e]r^N  (hh�eeee]r_N  (hheeejRN  jRN  jRN  jRN  ]r`N  (jYF  ]raN  (j[F  ]rbN  (j]F  ]rcN  (h	h�e]rdN  (hh�e]reN  (hhe]rfN  (jdF  ]rgN  (h	he]rhN  (hh�e]riN  (hhe]rjN  (j�K  ]rkN  (h	h�e]rlN  (hh�eeee]rmN  (hheeej`N  j`N  ]rnN  (jYF  ]roN  (j[F  ]rpN  (j]F  ]rqN  (h	h�e]rrN  (hh�e]rsN  (hhe]rtN  (jdF  ]ruN  (h	he]rvN  (hh�e]rwN  (hhe]rxN  (j�K  ]ryN  (h	h�e]rzN  (hh�eeee]r{N  (hheeejnN  jnN  jnN  jnN  ]r|N  (jYF  ]r}N  (j[F  ]r~N  (j]F  ]rN  (h	h�e]r�N  (hh�e]r�N  (hhe]r�N  (jdF  ]r�N  (h	he]r�N  (hh�e]r�N  (hhe]r�N  (j�K  ]r�N  (h	h�e]r�N  (hh�eeee]r�N  (hheee]r�N  (jYF  ]r�N  (j[F  ]r�N  (j]F  ]r�N  (h	h�e]r�N  (hh�e]r�N  (hhe]r�N  (jdF  ]r�N  (h	he]r�N  (hh�e]r�N  (hhe]r�N  (j�K  ]r�N  (h	h�e]r�N  (hh�eeee]r�N  (hheeej�N  j�N  j�N  ]r�N  (jYF  ]r�N  (j[F  ]r�N  (j]F  ]r�N  (h	j�  e]r�N  (hh�e]r�N  (hhe]r�N  (jdF  ]r�N  (h	he]r�N  (hh�e]r�N  (hhe]r�N  (j�K  ]r�N  (h	h�e]r�N  (hh�eeee]r�N  (hheeej�N  j�N  j�N  j�N  j�N  j�N  ]r�N  (jYF  ]r�N  (j[F  ]r�N  (j]F  ]r�N  (h	j�  e]r�N  (hh�e]r�N  (hhe]r�N  (jdF  ]r�N  (h	he]r�N  (hh�e]r�N  (hhe]r�N  (j�K  ]r�N  (h	h�e]r�N  (hh�eeee]r�N  (hheeej�N  j�N  j�N  j�N  j�N  ]r�N  (jYF  ]r�N  (j[F  ]r�N  (j]F  ]r�N  (h	j�  e]r�N  (hh�e]r�N  (hhe]r�N  (jdF  ]r�N  (h	he]r�N  (hh�e]r�N  (hhe]r�N  (j�K  ]r�N  (h	h�e]r�N  (hh�eeee]r�N  (hheeej�N  ]r�N  (jYF  ]r�N  (j[F  ]r�N  (j]F  ]r�N  (h	j�  e]r�N  (hh�e]r�N  (hhe]r�N  (jdF  ]r�N  (h	he]r�N  (hh�e]r�N  (hhe]r�N  (j�K  ]r�N  (h	h�e]r�N  (hh�eeee]r�N  (hheeej�N  j�N  j�N  j�N  j�N  j�N  j�N  ]r�N  (jYF  ]r�N  (j[F  ]r�N  (j]F  ]r�N  (h	j�  e]r�N  (hh�e]r�N  (hhe]r�N  (jdF  ]r�N  (h	he]r�N  (hh�e]r�N  (hhe]r�N  (j�K  ]r�N  (h	h�e]r�N  (hh�eeee]r�N  (hheeej�N  ]r�N  (jYF  ]r�N  (j[F  ]r�N  (j]F  ]r�N  (h	j�  e]r�N  (hh�e]r�N  (hhe]r�N  (jdF  ]r�N  (h	he]r�N  (hh�e]r�N  (hhe]r�N  (j�K  ]r�N  (h	h�e]r�N  (hh�eeee]r�N  (hheeej�N  j�N  ]r�N  (jYF  ]r�N  (j[F  ]r�N  (j]F  ]r�N  (h	j�  e]r�N  (hh�e]r�N  (hhe]r�N  (jdF  ]r�N  (h	he]r�N  (hh�e]r�N  (hhe]r�N  (j�K  ]r�N  (h	h�e]r�N  (hh�eeee]r�N  (hheeej�N  j�N  j�N  j�N  j�N  j�N  j�N  j�N  j�N  j�N  j�N  ]r�N  (jYF  ]r�N  (j[F  ]r�N  (j]F  ]r�N  (h	j�  e]r�N  (hh�e]r�N  (hhe]r O  (jdF  ]rO  (h	he]rO  (hh�e]rO  (hhe]rO  (j�K  ]rO  (h	h�e]rO  (hh�eeee]rO  (hheeej�N  j�N  j�N  ]rO  (jYF  ]r	O  (j[F  ]r
O  (j]F  ]rO  (h	j�  e]rO  (hh�e]rO  (hhe]rO  (jdF  ]rO  (h	he]rO  (hh�e]rO  (hhe]rO  (j�K  ]rO  (h	h�e]rO  (hh�eeee]rO  (hheeejO  ]rO  (jYF  ]rO  (j[F  ]rO  (j]F  ]rO  (h	j�  e]rO  (hh�e]rO  (hhe]rO  (jdF  ]rO  (h	he]rO  (hh�e]rO  (hhe]r O  (j�K  ]r!O  (h	h�e]r"O  (hh�eeee]r#O  (hheeejO  ]r$O  (jYF  ]r%O  (j[F  ]r&O  (j]F  ]r'O  (h	j�  e]r(O  (hh�e]r)O  (hhe]r*O  (jdF  ]r+O  (h	he]r,O  (hh�e]r-O  (hhe]r.O  (j�K  ]r/O  (h	h�e]r0O  (hh�eeee]r1O  (hheeej$O  j$O  j$O  j$O  j$O  j$O  j$O  j$O  j$O  ]r2O  (jYF  ]r3O  (j[F  ]r4O  (j]F  ]r5O  (h	j�  e]r6O  (hh�e]r7O  (hhe]r8O  (jdF  ]r9O  (h	he]r:O  (hh�e]r;O  (hhe]r<O  (j�K  ]r=O  (h	h�e]r>O  (hh�eeee]r?O  (hheeej2O  ]r@O  (jYF  ]rAO  (j[F  ]rBO  (j]F  ]rCO  (h	j�  e]rDO  (hh�e]rEO  (hhe]rFO  (jdF  ]rGO  (h	he]rHO  (hh�e]rIO  (hhe]rJO  (j�K  ]rKO  (h	h�e]rLO  (hh�eeee]rMO  (hheeej@O  j@O  j@O  j@O  ]rNO  (jYF  ]rOO  (j[F  ]rPO  (j]F  ]rQO  (h	j�  e]rRO  (hh�e]rSO  (hhe]rTO  (jdF  ]rUO  (h	he]rVO  (hh�e]rWO  (hhe]rXO  (j�K  ]rYO  (h	h�e]rZO  (hh�eeee]r[O  (hheeejNO  jNO  jNO  jNO  ]r\O  (jYF  ]r]O  (j[F  ]r^O  (j]F  ]r_O  (h	j�  e]r`O  (hh�e]raO  (hhe]rbO  (jdF  ]rcO  (h	he]rdO  (hh�e]reO  (hhe]rfO  (j�K  ]rgO  (h	h�e]rhO  (hh�eeee]riO  (hheeej\O  j\O  ]rjO  (jYF  ]rkO  (j[F  ]rlO  (j]F  ]rmO  (h	j�  e]rnO  (hh�e]roO  (hhe]rpO  (jdF  ]rqO  (h	he]rrO  (hh�e]rsO  (hhe]rtO  (j�K  ]ruO  (h	h�e]rvO  (hh�eeee]rwO  (hheeejjO  jjO  jjO  ]rxO  (jYF  ]ryO  (j[F  ]rzO  (j]F  ]r{O  (h	j�  e]r|O  (hh�e]r}O  (hhe]r~O  (jdF  ]rO  (h	he]r�O  (hh�e]r�O  (hhe]r�O  (j�K  ]r�O  (h	h�e]r�O  (hh�eeee]r�O  (hheeejxO  ]r�O  (jYF  ]r�O  (j[F  ]r�O  (j]F  ]r�O  (h	j�  e]r�O  (hh�e]r�O  (hhe]r�O  (jdF  ]r�O  (h	he]r�O  (hh�e]r�O  (hhe]r�O  (j�K  ]r�O  (h	h�e]r�O  (hh�eeee]r�O  (hheeej�O  j�O  j�O  j�O  j�O  j�O  ]r�O  (jYF  ]r�O  (j[F  ]r�O  (j]F  ]r�O  (h	j�  e]r�O  (hh�e]r�O  (hhe]r�O  (jdF  ]r�O  (h	he]r�O  (hh�e]r�O  (hhe]r�O  (j�K  ]r�O  (h	h�e]r�O  (hh�eeee]r�O  (hheee]r�O  (jYF  ]r�O  (j[F  ]r�O  (j]F  ]r�O  (h	j�  e]r�O  (hh�e]r�O  (hhe]r�O  (jdF  ]r�O  (h	he]r�O  (hh�e]r�O  (hhe]r�O  (j�K  ]r�O  (h	h�e]r�O  (hh�eeee]r�O  (hheeej�O  j�O  j�O  j�O  j�O  j�O  j�O  ]r�O  (jYF  ]r�O  (j[F  ]r�O  (j]F  ]r�O  (h	j�  e]r�O  (hh�e]r�O  (hhe]r�O  (jdF  ]r�O  (h	he]r�O  (hh�e]r�O  (hhe]r�O  (j�K  ]r�O  (h	h�e]r�O  (hh�eeee]r�O  (hheeej�O  j�O  ]r�O  (jYF  ]r�O  (j[F  ]r�O  (j]F  ]r�O  (h	j�  e]r�O  (hh�e]r�O  (hhe]r�O  (jdF  ]r�O  (h	he]r�O  (hh�e]r�O  (hhe]r�O  (j�K  ]r�O  (h	h�e]r�O  (hh�eeee]r�O  (hheeej�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  ]r�O  (jYF  ]r�O  (j[F  ]r�O  (j]F  ]r�O  (h	j�  e]r�O  (hh�e]r�O  (hhe]r�O  (jdF  ]r�O  (h	he]r�O  (hh�e]r�O  (hhe]r�O  (j�K  ]r�O  (h	h�e]r�O  (hh�eeee]r�O  (hheeej�O  j�O  ]r�O  (jYF  ]r�O  (j[F  ]r�O  (j]F  ]r�O  (h	j�  e]r�O  (hh�e]r�O  (hhe]r�O  (jdF  ]r�O  (h	he]r�O  (hh�e]r�O  (hhe]r�O  (j�K  ]r�O  (h	h�e]r�O  (hh�eeee]r�O  (hheee]r�O  (jYF  ]r�O  (j[F  ]r�O  (j]F  ]r�O  (h	j�  e]r�O  (hh�e]r�O  (hhe]r�O  (jdF  ]r�O  (h	he]r�O  (hh�e]r�O  (hhe]r�O  (j�K  ]r�O  (h	h�e]r�O  (hh�eeee]r�O  (hheee]r�O  (jYF  ]r�O  (j[F  ]r�O  (j]F  ]r�O  (h	j�  e]r�O  (hh�e]r�O  (hhe]r�O  (jdF  ]r�O  (h	he]r�O  (hh�e]r�O  (hhe]r P  (j�K  ]rP  (h	h�e]rP  (hh�eeee]rP  (hheeej�O  j�O  ]rP  (jYF  ]rP  (j[F  ]rP  (j]F  ]rP  (h	j�  e]rP  (hh�e]r	P  (hhe]r
P  (jdF  ]rP  (h	he]rP  (hh�e]rP  (hhe]rP  (j�K  ]rP  (h	h�e]rP  (hh�eeee]rP  (hheee]rP  (jYF  ]rP  (j[F  ]rP  (j]F  ]rP  (h	j�  e]rP  (hh�e]rP  (hhe]rP  (jdF  ]rP  (h	he]rP  (hh�e]rP  (hhe]rP  (j�K  ]rP  (h	h�e]rP  (hh�eeee]rP  (hheeejP  jP  jP  jP  jP  ]r P  (jYF  ]r!P  (j[F  ]r"P  (j]F  ]r#P  (h	j�  e]r$P  (hh�e]r%P  (hhe]r&P  (jdF  ]r'P  (h	he]r(P  (hh�e]r)P  (hhe]r*P  (j�K  ]r+P  (h	h�e]r,P  (hh�eeee]r-P  (hheeej P  ]r.P  (jYF  ]r/P  (j[F  ]r0P  (j]F  ]r1P  (h	j�  e]r2P  (hh�e]r3P  (hhe]r4P  (jdF  ]r5P  (h	he]r6P  (hh�e]r7P  (hhe]r8P  (j�K  ]r9P  (h	h�e]r:P  (hh�eeee]r;P  (hheeej.P  ]r<P  (jYF  ]r=P  (j[F  ]r>P  (j]F  ]r?P  (h	j�  e]r@P  (hh�e]rAP  (hhe]rBP  (jdF  ]rCP  (h	he]rDP  (hh�e]rEP  (hhe]rFP  (j�K  ]rGP  (h	h�e]rHP  (hh�eeee]rIP  (hheeej<P  j<P  j<P  j<P  ]rJP  (jYF  ]rKP  (j[F  ]rLP  (j]F  ]rMP  (h	j�  e]rNP  (hh�e]rOP  (hhe]rPP  (jdF  ]rQP  (h	he]rRP  (hh�e]rSP  (hhe]rTP  (j�K  ]rUP  (h	h�e]rVP  (hh�eeee]rWP  (hheeejJP  ]rXP  (jYF  ]rYP  (j[F  ]rZP  (j]F  ]r[P  (h	h�e]r\P  (hh�e]r]P  (hhe]r^P  (jdF  ]r_P  (h	he]r`P  (hh�e]raP  (hhe]rbP  (j�K  ]rcP  (h	h�e]rdP  (hh�eeee]reP  (hheeejXP  jXP  jXP  ]rfP  (jYF  ]rgP  (j[F  ]rhP  (j]F  ]riP  (h	h�e]rjP  (hh�e]rkP  (hhe]rlP  (jdF  ]rmP  (h	he]rnP  (hh�e]roP  (hhe]rpP  (j�K  ]rqP  (h	h�e]rrP  (hh�eeee]rsP  (hheee]rtP  (jYF  ]ruP  (j[F  ]rvP  (j]F  ]rwP  (h	j�  e]rxP  (hh�e]ryP  (hhe]rzP  (jdF  ]r{P  (h	he]r|P  (hh�e]r}P  (hhe]r~P  (j�K  ]rP  (h	h�e]r�P  (hh�eeee]r�P  (hheeejtP  jtP  jtP  ]r�P  (jYF  ]r�P  (j[F  ]r�P  (j]F  ]r�P  (h	j�  e]r�P  (hh�e]r�P  (hhe]r�P  (jdF  ]r�P  (h	he]r�P  (hh�e]r�P  (hhe]r�P  (j�K  ]r�P  (h	h�e]r�P  (hh�eeee]r�P  (hheeej�P  j�P  ]r�P  (jYF  ]r�P  (j[F  ]r�P  (j]F  ]r�P  (h	j�  e]r�P  (hh�e]r�P  (hhe]r�P  (jdF  ]r�P  (h	he]r�P  (hh�e]r�P  (hhe]r�P  (j�K  ]r�P  (h	h�e]r�P  (hh�eeee]r�P  (hheeej�P  j�P  j�P  ]r�P  (jYF  ]r�P  (j[F  ]r�P  (j]F  ]r�P  (h	j�  e]r�P  (hh�e]r�P  (hhe]r�P  (jdF  ]r�P  (h	he]r�P  (hh�e]r�P  (hhe]r�P  (j�K  ]r�P  (h	h�e]r�P  (hh�eeee]r�P  (hheeej�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  ]r�P  (jYF  ]r�P  (j[F  ]r�P  (j]F  ]r�P  (h	j�  e]r�P  (hh�e]r�P  (hhe]r�P  (jdF  ]r�P  (h	he]r�P  (hh�e]r�P  (hhe]r�P  (j�K  ]r�P  (h	h�e]r�P  (hh�eeee]r�P  (hheeej�P  j�P  ]r�P  (jYF  ]r�P  (j[F  ]r�P  (j]F  ]r�P  (h	j�  e]r�P  (hh�e]r�P  (hhe]r�P  (jdF  ]r�P  (h	he]r�P  (hh�e]r�P  (hhe]r�P  (j�K  ]r�P  (h	h�e]r�P  (hh�eeee]r�P  (hheeej�P  j�P  j�P  j�P  j�P  ]r�P  (jYF  ]r�P  (j[F  ]r�P  (j]F  ]r�P  (h	j�  e]r�P  (hh�e]r�P  (hhe]r�P  (jdF  ]r�P  (h	he]r�P  (hh�e]r�P  (hhe]r�P  (j�K  ]r�P  (h	h�e]r�P  (hh�eeee]r�P  (hheee]r�P  (jYF  ]r�P  (j[F  ]r�P  (j]F  ]r�P  (h	j�  e]r�P  (hh�e]r�P  (hhe]r�P  (jdF  ]r�P  (h	he]r�P  (hh�e]r�P  (hhe]r�P  (j�K  ]r�P  (h	h�e]r�P  (hh�eeee]r�P  (hheee]r�P  (jYF  ]r�P  (j[F  ]r�P  (j]F  ]r�P  (h	j�  e]r�P  (hh�e]r�P  (hhe]r�P  (jdF  ]r�P  (h	he]r�P  (hh�e]r�P  (hhe]r�P  (j�K  ]r�P  (h	h�e]r�P  (hh�eeee]r�P  (hheee]r�P  (jYF  ]r�P  (j[F  ]r�P  (j]F  ]r�P  (h	j�  e]r�P  (hh�e]r�P  (hhe]r�P  (jdF  ]r�P  (h	he]r�P  (hh�e]r�P  (hhe]r�P  (j�K  ]r�P  (h	h�e]r�P  (hh�eeee]r�P  (hheeej�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  j�P  ]r Q  (jYF  ]rQ  (j[F  ]rQ  (j]F  ]rQ  (h	j�  e]rQ  (hh�e]rQ  (hhe]rQ  (jdF  ]rQ  (h	he]rQ  (hh�e]r	Q  (hhe]r
Q  (j�K  ]rQ  (h	h�e]rQ  (hh�eeee]rQ  (hheeej Q  j Q  j Q  j Q  j Q  j Q  j Q  j Q  j Q  j Q  j Q  j Q  j Q  j Q  j Q  j Q  j Q  j Q  ]rQ  (jYF  ]rQ  (j[F  ]rQ  (j]F  ]rQ  (h	j�  e]rQ  (hh�e]rQ  (hhe]rQ  (jdF  ]rQ  (h	he]rQ  (hh�e]rQ  (hhe]rQ  (j�K  ]rQ  (h	h�e]rQ  (hh�eeee]rQ  (hheeejQ  jQ  jQ  jQ  jQ  ]rQ  (jYF  ]rQ  (j[F  ]rQ  (j]F  ]rQ  (h	j�  e]r Q  (hh�e]r!Q  (hhe]r"Q  (jdF  ]r#Q  (h	he]r$Q  (hh�e]r%Q  (hhe]r&Q  (j�K  ]r'Q  (h	h�e]r(Q  (hh�eeee]r)Q  (hheeejQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  ]r*Q  (jYF  ]r+Q  (j[F  ]r,Q  (j]F  ]r-Q  (h	j�  e]r.Q  (hh�e]r/Q  (hhe]r0Q  (jdF  ]r1Q  (h	he]r2Q  (hh�e]r3Q  (hhe]r4Q  (j�K  ]r5Q  (h	h�e]r6Q  (hh�eeee]r7Q  (hheeej*Q  j*Q  j*Q  ]r8Q  (jYF  ]r9Q  (j[F  ]r:Q  (j]F  ]r;Q  (h	j�  e]r<Q  (hh�e]r=Q  (hhe]r>Q  (jdF  ]r?Q  (h	he]r@Q  (hh�e]rAQ  (hhe]rBQ  (j�K  ]rCQ  (h	h�e]rDQ  (hh�eeee]rEQ  (hheeej8Q  j8Q  ]rFQ  (jYF  ]rGQ  (j[F  ]rHQ  (j]F  ]rIQ  (h	j�  e]rJQ  (hh�e]rKQ  (hhe]rLQ  (jdF  ]rMQ  (h	he]rNQ  (hh�e]rOQ  (hhe]rPQ  (j�K  ]rQQ  (h	h�e]rRQ  (hh�eeee]rSQ  (hheeejFQ  jFQ  jFQ  jFQ  jFQ  jFQ  jFQ  ]rTQ  (jYF  ]rUQ  (j[F  ]rVQ  (j]F  ]rWQ  (h	j�  e]rXQ  (hh�e]rYQ  (hhe]rZQ  (jdF  ]r[Q  (h	he]r\Q  (hh�e]r]Q  (hhe]r^Q  (j�K  ]r_Q  (h	h�e]r`Q  (hh�eeee]raQ  (hheee]rbQ  (jYF  ]rcQ  (j[F  ]rdQ  (j]F  ]reQ  (h	j�  e]rfQ  (hh�e]rgQ  (hhe]rhQ  (jdF  ]riQ  (h	he]rjQ  (hh�e]rkQ  (hhe]rlQ  (X	   Next-MovermQ  ]rnQ  (h	h�e]roQ  (hh�eeee]rpQ  (hheeejbQ  jbQ  jbQ  jbQ  jbQ  jbQ  jbQ  jbQ  jbQ  jbQ  jbQ  jbQ  jbQ  jbQ  jbQ  jbQ  ]rqQ  (jYF  ]rrQ  (j[F  ]rsQ  (j]F  ]rtQ  (h	j�  e]ruQ  (hh�e]rvQ  (hhe]rwQ  (jdF  ]rxQ  (h	he]ryQ  (hh�e]rzQ  (hhe]r{Q  (jmQ  ]r|Q  (h	h�e]r}Q  (hh�eeee]r~Q  (hheee]rQ  (jYF  ]r�Q  (j[F  ]r�Q  (j]F  ]r�Q  (h	j�  e]r�Q  (hh�e]r�Q  (hhe]r�Q  (jdF  ]r�Q  (h	he]r�Q  (hh�e]r�Q  (hhe]r�Q  (jmQ  ]r�Q  (h	h�e]r�Q  (hh�eeee]r�Q  (hheeejQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  jQ  ]r�Q  (jYF  ]r�Q  (j[F  ]r�Q  (j]F  ]r�Q  (h	j�  e]r�Q  (hh�e]r�Q  (hhe]r�Q  (jdF  ]r�Q  (h	he]r�Q  (hh�e]r�Q  (hhe]r�Q  (jmQ  ]r�Q  (h	h�e]r�Q  (hh�eeee]r�Q  (hheeej�Q  ]r�Q  (jYF  ]r�Q  (j[F  ]r�Q  (j]F  ]r�Q  (h	j�  e]r�Q  (hh�e]r�Q  (hhe]r�Q  (jdF  ]r�Q  (h	he]r�Q  (hh�e]r�Q  (hhe]r�Q  (jmQ  ]r�Q  (h	h�e]r�Q  (hh�eeee]r�Q  (hheeej�Q  j�Q  j�Q  j�Q  j�Q  ]r�Q  (jYF  ]r�Q  (j[F  ]r�Q  (j]F  ]r�Q  (h	j�  e]r�Q  (hh�e]r�Q  (hhe]r�Q  (jdF  ]r�Q  (h	he]r�Q  (hh�e]r�Q  (hhe]r�Q  (jmQ  ]r�Q  (h	h�e]r�Q  (hh�eeee]r�Q  (hheeej�Q  j�Q  j�Q  j�Q  j�Q  j�Q  j�Q  ]r�Q  (jYF  ]r�Q  (j[F  ]r�Q  (j]F  ]r�Q  (h	j�  e]r�Q  (hh�e]r�Q  (hhe]r�Q  (jdF  ]r�Q  (h	he]r�Q  (hh�e]r�Q  (hhe]r�Q  (jmQ  ]r�Q  (h	h�e]r�Q  (hh�eeee]r�Q  (hheeej�Q  j�Q  j�Q  ]r�Q  (jYF  ]r�Q  (j[F  ]r�Q  (j]F  ]r�Q  (h	j�  e]r�Q  (hh�e]r�Q  (hhe]r�Q  (jdF  ]r�Q  (h	he]r�Q  (hh�e]r�Q  (hhe]r�Q  (jmQ  ]r�Q  (h	h�e]r�Q  (hh�eeee]r�Q  (hheee]r�Q  (jYF  ]r�Q  (j[F  ]r�Q  (j]F  ]r�Q  (h	j�  e]r�Q  (hh�e]r�Q  (hhe]r�Q  (jdF  ]r�Q  (h	he]r�Q  (hh�e]r�Q  (hhe]r�Q  (jmQ  ]r�Q  (h	h�e]r�Q  (hh�eeee]r�Q  (hheeej�Q  j�Q  ]r�Q  (jYF  ]r�Q  (j[F  ]r�Q  (j]F  ]r�Q  (h	j�  e]r�Q  (hh�e]r�Q  (hhe]r�Q  (jdF  ]r�Q  (h	he]r�Q  (hh�e]r�Q  (hhe]r�Q  (jmQ  ]r�Q  (h	h�e]r�Q  (hh�eeee]r�Q  (hheeej�Q  j�Q  j�Q  j�Q  j�Q  j�Q  j�Q  j�Q  ]r�Q  (jYF  ]r�Q  (j[F  ]r�Q  (j]F  ]r�Q  (h	j�  e]r�Q  (hh�e]r�Q  (hhe]r�Q  (jdF  ]r�Q  (h	he]r�Q  (hh�e]r�Q  (hhe]r�Q  (jmQ  ]r�Q  (h	h�e]r�Q  (hh�eeee]r�Q  (hheeej�Q  j�Q  j�Q  j�Q  j�Q  j�Q  j�Q  ]r�Q  (jYF  ]r�Q  (j[F  ]r�Q  (j]F  ]r R  (h	j�  e]rR  (hh�e]rR  (hhe]rR  (jdF  ]rR  (h	he]rR  (hh�e]rR  (hhe]rR  (jmQ  ]rR  (h	h�e]r	R  (hh�eeee]r
R  (hheeej�Q  j�Q  j�Q  ]rR  (jYF  ]rR  (j[F  ]rR  (j]F  ]rR  (h	j�  e]rR  (hh�e]rR  (hhe]rR  (jdF  ]rR  (h	he]rR  (hh�e]rR  (hhe]rR  (jmQ  ]rR  (h	h�e]rR  (hh�eeee]rR  (hheeejR  jR  jR  jR  jR  ]rR  (jYF  ]rR  (j[F  ]rR  (j]F  ]rR  (h	j�  e]rR  (hh�e]rR  (hhe]rR  (jdF  ]r R  (h	he]r!R  (hh�e]r"R  (hhe]r#R  (jmQ  ]r$R  (h	h�e]r%R  (hh�eeee]r&R  (hheee]r'R  (jYF  ]r(R  (j[F  ]r)R  (j]F  ]r*R  (h	j�  e]r+R  (hh�e]r,R  (hhe]r-R  (jdF  ]r.R  (h	he]r/R  (hh�e]r0R  (hhe]r1R  (X	   Next-Mover2R  ]r3R  (h	h�e]r4R  (hh�eeee]r5R  (hheeej'R  j'R  j'R  j'R  j'R  j'R  ]r6R  (jYF  ]r7R  (j[F  ]r8R  (j]F  ]r9R  (h	j�  e]r:R  (hh�e]r;R  (hhe]r<R  (jdF  ]r=R  (h	he]r>R  (hh�e]r?R  (hhe]r@R  (j2R  ]rAR  (h	h�e]rBR  (hh�eeee]rCR  (hheee]rDR  (jYF  ]rER  (j[F  ]rFR  (j]F  ]rGR  (h	j�  e]rHR  (hh�e]rIR  (hhe]rJR  (jdF  ]rKR  (h	he]rLR  (hh�e]rMR  (hhe]rNR  (j2R  ]rOR  (h	h�e]rPR  (hh�eeee]rQR  (hheeejDR  ]rRR  (jYF  ]rSR  (j[F  ]rTR  (j]F  ]rUR  (h	j�  e]rVR  (hh�e]rWR  (hhe]rXR  (jdF  ]rYR  (h	he]rZR  (hh�e]r[R  (hhe]r\R  (j2R  ]r]R  (h	h�e]r^R  (hh�eeee]r_R  (hheee]r`R  (jYF  ]raR  (j[F  ]rbR  (j]F  ]rcR  (h	j�  e]rdR  (hh�e]reR  (hhe]rfR  (jdF  ]rgR  (h	he]rhR  (hh�e]riR  (hhe]rjR  (j2R  ]rkR  (h	h�e]rlR  (hh�eeee]rmR  (hheeej`R  ]rnR  (jYF  ]roR  (j[F  ]rpR  (j]F  ]rqR  (h	j�  e]rrR  (hh�e]rsR  (hhe]rtR  (jdF  ]ruR  (h	he]rvR  (hh�e]rwR  (hhe]rxR  (j2R  ]ryR  (h	h�e]rzR  (hh�eeee]r{R  (hheee]r|R  (jYF  ]r}R  (j[F  ]r~R  (j]F  ]rR  (h	j�  e]r�R  (hh�e]r�R  (hhe]r�R  (jdF  ]r�R  (h	he]r�R  (hh�e]r�R  (hhe]r�R  (j2R  ]r�R  (h	h�e]r�R  (hh�eeee]r�R  (hheee]r�R  (jYF  ]r�R  (j[F  ]r�R  (j]F  ]r�R  (h	j�  e]r�R  (hh�e]r�R  (hhe]r�R  (jdF  ]r�R  (h	he]r�R  (hh�e]r�R  (hhe]r�R  (j2R  ]r�R  (h	h�e]r�R  (hh�eeee]r�R  (hheeej�R  j�R  j�R  j�R  j�R  j�R  j�R  j�R  j�R  j�R  j�R  ]r�R  (jYF  ]r�R  (j[F  ]r�R  (j]F  ]r�R  (h	j�  e]r�R  (hh�e]r�R  (hhe]r�R  (jdF  ]r�R  (h	he]r�R  (hh�e]r�R  (hhe]r�R  (j2R  ]r�R  (h	h�e]r�R  (hh�eeee]r�R  (hheeej�R  j�R  j�R  j�R  j�R  j�R  j�R  j�R  ]r�R  (jYF  ]r�R  (j[F  ]r�R  (j]F  ]r�R  (h	j�  e]r�R  (hh�e]r�R  (hhe]r�R  (jdF  ]r�R  (h	he]r�R  (hh�e]r�R  (hhe]r�R  (j2R  ]r�R  (h	h�e]r�R  (hh�eeee]r�R  (hheeej�R  j�R  j�R  j�R  j�R  e(]r�R  (jYF  ]r�R  (j[F  ]r�R  (j]F  ]r�R  (h	j�  e]r�R  (hh�e]r�R  (hhe]r�R  (jdF  ]r�R  (h	he]r�R  (hh�e]r�R  (hhe]r�R  (j2R  ]r�R  (h	h�e]r�R  (hh�eeee]r�R  (hheee]r�R  (jYF  ]r�R  (j[F  ]r�R  (j]F  ]r�R  (h	j�  e]r�R  (hh�e]r�R  (hhe]r�R  (jdF  ]r�R  (h	he]r�R  (hh�e]r�R  (hhe]r�R  (j2R  ]r�R  (h	h�e]r�R  (hh�eeee]r�R  (hheeej�R  ]r�R  (jYF  ]r�R  (j[F  ]r�R  (j]F  ]r�R  (h	j�  e]r�R  (hh�e]r�R  (hhe]r�R  (jdF  ]r�R  (h	he]r�R  (hh�e]r�R  (hhe]r�R  (j2R  ]r�R  (h	h�e]r�R  (hh�eeee]r�R  (hheee]r�R  (jYF  ]r�R  (j[F  ]r�R  (j]F  ]r�R  (h	j�  e]r�R  (hh�e]r�R  (hhe]r�R  (jdF  ]r�R  (h	he]r�R  (hh�e]r�R  (hhe]r�R  (j2R  ]r�R  (h	h�e]r�R  (hh�eeee]r�R  (hheeej�R  j�R  ]r�R  (jYF  ]r�R  (j[F  ]r�R  (j]F  ]r�R  (h	j�  e]r�R  (hh�e]r�R  (hhe]r�R  (jdF  ]r�R  (h	he]r�R  (hh�e]r�R  (hhe]r�R  (j2R  ]r�R  (h	h�e]r�R  (hh�eeee]r�R  (hheee]r�R  (jYF  ]r�R  (j[F  ]r�R  (j]F  ]r�R  (h	j�  e]r�R  (hh�e]r�R  (hhe]r S  (jdF  ]rS  (h	he]rS  (hh�e]rS  (hhe]rS  (j2R  ]rS  (h	h�e]rS  (hh�eeee]rS  (hheee]rS  (jYF  ]r	S  (j[F  ]r
S  (j]F  ]rS  (h	j�  e]rS  (hh�e]rS  (hhe]rS  (jdF  ]rS  (h	he]rS  (hh�e]rS  (hhe]rS  (j2R  ]rS  (h	h�e]rS  (hh�eeee]rS  (hheee]rS  (jYF  ]rS  (j[F  ]rS  (j]F  ]rS  (h	j�  e]rS  (hh�e]rS  (hhe]rS  (jdF  ]rS  (h	he]rS  (hh�e]rS  (hhe]r S  (j2R  ]r!S  (h	h�e]r"S  (hh�eeee]r#S  (hheeejS  jS  jS  ]r$S  (jYF  ]r%S  (j[F  ]r&S  (j]F  ]r'S  (h	j�  e]r(S  (hh�e]r)S  (hhe]r*S  (jdF  ]r+S  (h	he]r,S  (hh�e]r-S  (hhe]r.S  (j2R  ]r/S  (h	h�e]r0S  (hh�eeee]r1S  (hheeej$S  j$S  j$S  j$S  j$S  j$S  j$S  j$S  ]r2S  (jYF  ]r3S  (j[F  ]r4S  (j]F  ]r5S  (h	j�  e]r6S  (hh�e]r7S  (hhe]r8S  (jdF  ]r9S  (h	he]r:S  (hh�e]r;S  (hhe]r<S  (j2R  ]r=S  (h	h�e]r>S  (hh�eeee]r?S  (hheeej2S  j2S  j2S  ]r@S  (jYF  ]rAS  (j[F  ]rBS  (j]F  ]rCS  (h	j�  e]rDS  (hh�e]rES  (hhe]rFS  (jdF  ]rGS  (h	he]rHS  (hh�e]rIS  (hhe]rJS  (j2R  ]rKS  (h	h�e]rLS  (hh�eeee]rMS  (hheeej@S  j@S  j@S  j@S  j@S  j@S  ]rNS  (jYF  ]rOS  (j[F  ]rPS  (j]F  ]rQS  (h	j�  e]rRS  (hh�e]rSS  (hhe]rTS  (jdF  ]rUS  (h	he]rVS  (hh�e]rWS  (hhe]rXS  (j2R  ]rYS  (h	h�e]rZS  (hh�eeee]r[S  (hheeejNS  jNS  jNS  jNS  jNS  ]r\S  (jYF  ]r]S  (j[F  ]r^S  (j]F  ]r_S  (h	j�  e]r`S  (hh�e]raS  (hhe]rbS  (jdF  ]rcS  (h	he]rdS  (hh�e]reS  (hhe]rfS  (j2R  ]rgS  (h	h�e]rhS  (hh�eeee]riS  (hheee]rjS  (jYF  ]rkS  (j[F  ]rlS  (j]F  ]rmS  (h	j�  e]rnS  (hh�e]roS  (hhe]rpS  (jdF  ]rqS  (h	he]rrS  (hh�e]rsS  (hhe]rtS  (j2R  ]ruS  (h	h�e]rvS  (hh�eeee]rwS  (hheee]rxS  (jYF  ]ryS  (j[F  ]rzS  (j]F  ]r{S  (h	j�  e]r|S  (hh�e]r}S  (hhe]r~S  (jdF  ]rS  (h	he]r�S  (hh�e]r�S  (hhe]r�S  (j2R  ]r�S  (h	h�e]r�S  (hh�eeee]r�S  (hheee]r�S  (jYF  ]r�S  (j[F  ]r�S  (j]F  ]r�S  (h	j�  e]r�S  (hh�e]r�S  (hhe]r�S  (jdF  ]r�S  (h	he]r�S  (hh�e]r�S  (hhe]r�S  (j2R  ]r�S  (h	h�e]r�S  (hh�eeee]r�S  (hheeej�S  j�S  j�S  ]r�S  (jYF  ]r�S  (j[F  ]r�S  (j]F  ]r�S  (h	j�  e]r�S  (hh�e]r�S  (hhe]r�S  (jdF  ]r�S  (h	he]r�S  (hh�e]r�S  (hhe]r�S  (j2R  ]r�S  (h	h�e]r�S  (hh�eeee]r�S  (hheee]r�S  (jYF  ]r�S  (j[F  ]r�S  (j]F  ]r�S  (h	j�  e]r�S  (hh�e]r�S  (hhe]r�S  (jdF  ]r�S  (h	he]r�S  (hh�e]r�S  (hhe]r�S  (j2R  ]r�S  (h	h�e]r�S  (hh�eeee]r�S  (hheee]r�S  (jYF  ]r�S  (j[F  ]r�S  (j]F  ]r�S  (h	j�  e]r�S  (hh�e]r�S  (hhe]r�S  (jdF  ]r�S  (h	he]r�S  (hh�e]r�S  (hhe]r�S  (j2R  ]r�S  (h	h�e]r�S  (hh�eeee]r�S  (hheeej�S  j�S  j�S  ]r�S  (jYF  ]r�S  (j[F  ]r�S  (j]F  ]r�S  (h	j�  e]r�S  (hh�e]r�S  (hhe]r�S  (jdF  ]r�S  (h	he]r�S  (hh�e]r�S  (hhe]r�S  (j2R  ]r�S  (h	h�e]r�S  (hh�eeee]r�S  (hheeej�S  j�S  j�S  j�S  j�S  j�S  j�S  j�S  j�S  j�S  j�S  j�S  j�S  ]r�S  (jYF  ]r�S  (j[F  ]r�S  (j]F  ]r�S  (h	j�  e]r�S  (hh�e]r�S  (hhe]r�S  (jdF  ]r�S  (h	he]r�S  (hh�e]r�S  (hhe]r�S  (j2R  ]r�S  (h	h�e]r�S  (hh�eeee]r�S  (hheee]r�S  (jYF  ]r�S  (j[F  ]r�S  (j]F  ]r�S  (h	j�  e]r�S  (hh�e]r�S  (hhe]r�S  (jdF  ]r�S  (h	he]r�S  (hh�e]r�S  (hhe]r�S  (j2R  ]r�S  (h	h�e]r�S  (hh�eeee]r�S  (hheeej�S  j�S  ]r�S  (jYF  ]r�S  (j[F  ]r�S  (j]F  ]r�S  (h	j�  e]r�S  (hh�e]r�S  (hhe]r�S  (jdF  ]r�S  (h	he]r�S  (hh�e]r�S  (hhe]r�S  (j2R  ]r�S  (h	h�e]r�S  (hh�eeee]r�S  (hheeej�S  j�S  j�S  ]r�S  (jYF  ]r�S  (j[F  ]r�S  (j]F  ]r�S  (h	j�  e]r�S  (hh�e]r�S  (hhe]r�S  (jdF  ]r�S  (h	he]r�S  (hh�e]r�S  (hhe]r T  (j2R  ]rT  (h	h�e]rT  (hh�eeee]rT  (hheeej�S  j�S  j�S  j�S  j�S  j�S  j�S  j�S  j�S  ]rT  (jYF  ]rT  (j[F  ]rT  (j]F  ]rT  (h	j�  e]rT  (hh�e]r	T  (hhe]r
T  (jdF  ]rT  (h	he]rT  (hh�e]rT  (hhe]rT  (j2R  ]rT  (h	h�e]rT  (hh�eeee]rT  (hheee]rT  (jYF  ]rT  (j[F  ]rT  (j]F  ]rT  (h	j�  e]rT  (hh�e]rT  (hhe]rT  (jdF  ]rT  (h	he]rT  (hh�e]rT  (hhe]rT  (j2R  ]rT  (h	h�e]rT  (hh�eeee]rT  (hheeejT  jT  jT  jT  ]r T  (jYF  ]r!T  (j[F  ]r"T  (j]F  ]r#T  (h	j�  e]r$T  (hh�e]r%T  (hhe]r&T  (jdF  ]r'T  (h	he]r(T  (hh�e]r)T  (hhe]r*T  (j2R  ]r+T  (h	h�e]r,T  (hh�eeee]r-T  (hheee]r.T  (jYF  ]r/T  (j[F  ]r0T  (j]F  ]r1T  (h	j�  e]r2T  (hh�e]r3T  (hhe]r4T  (jdF  ]r5T  (h	he]r6T  (hh�e]r7T  (hhe]r8T  (j2R  ]r9T  (h	h�e]r:T  (hh�eeee]r;T  (hheeej.T  ]r<T  (jYF  ]r=T  (j[F  ]r>T  (j]F  ]r?T  (h	j�  e]r@T  (hh�e]rAT  (hhe]rBT  (jdF  ]rCT  (h	he]rDT  (hh�e]rET  (hhe]rFT  (j2R  ]rGT  (h	h�e]rHT  (hh�eeee]rIT  (hheeej<T  j<T  j<T  j<T  j<T  j<T  j<T  j<T  j<T  j<T  j<T  ]rJT  (jYF  ]rKT  (j[F  ]rLT  (j]F  ]rMT  (h	j�  e]rNT  (hh�e]rOT  (hhe]rPT  (jdF  ]rQT  (h	he]rRT  (hh�e]rST  (hhe]rTT  (j2R  ]rUT  (h	h�e]rVT  (hh�eeee]rWT  (hheee]rXT  (jYF  ]rYT  (j[F  ]rZT  (j]F  ]r[T  (h	j�  e]r\T  (hh�e]r]T  (hhe]r^T  (jdF  ]r_T  (h	he]r`T  (hh�e]raT  (hhe]rbT  (j2R  ]rcT  (h	h�e]rdT  (hh�eeee]reT  (hheeejXT  ]rfT  (jYF  ]rgT  (j[F  ]rhT  (j]F  ]riT  (h	j�  e]rjT  (hh�e]rkT  (hhe]rlT  (jdF  ]rmT  (h	he]rnT  (hh�e]roT  (hhe]rpT  (j2R  ]rqT  (h	h�e]rrT  (hh�eeee]rsT  (hheeejfT  jfT  jfT  jfT  ]rtT  (jYF  ]ruT  (j[F  ]rvT  (j]F  ]rwT  (h	j�  e]rxT  (hh�e]ryT  (hhe]rzT  (jdF  ]r{T  (h	he]r|T  (hh�e]r}T  (hhe]r~T  (j2R  ]rT  (h	h�e]r�T  (hh�eeee]r�T  (hheeejtT  jtT  ]r�T  (jYF  ]r�T  (j[F  ]r�T  (j]F  ]r�T  (h	j�  e]r�T  (hh�e]r�T  (hhe]r�T  (jdF  ]r�T  (h	he]r�T  (hh�e]r�T  (hhe]r�T  (j2R  ]r�T  (h	h�e]r�T  (hh�eeee]r�T  (hheee]r�T  (jYF  ]r�T  (j[F  ]r�T  (j]F  ]r�T  (h	j�  e]r�T  (hh�e]r�T  (hhe]r�T  (jdF  ]r�T  (h	he]r�T  (hh�e]r�T  (hhe]r�T  (j2R  ]r�T  (h	h�e]r�T  (hh�eeee]r�T  (hheee]r�T  (jYF  ]r�T  (j[F  ]r�T  (j]F  ]r�T  (h	j�  e]r�T  (hh�e]r�T  (hhe]r�T  (jdF  ]r�T  (h	he]r�T  (hh�e]r�T  (hhe]r�T  (j2R  ]r�T  (h	h�e]r�T  (hh�eeee]r�T  (hheeej�T  j�T  j�T  ]r�T  (jYF  ]r�T  (j[F  ]r�T  (j]F  ]r�T  (h	j�  e]r�T  (hh�e]r�T  (hhe]r�T  (jdF  ]r�T  (h	he]r�T  (hh�e]r�T  (hhe]r�T  (j2R  ]r�T  (h	h�e]r�T  (hh�eeee]r�T  (hheee]r�T  (jYF  ]r�T  (j[F  ]r�T  (j]F  ]r�T  (h	j�  e]r�T  (hh�e]r�T  (hhe]r�T  (jdF  ]r�T  (h	he]r�T  (hh�e]r�T  (hhe]r�T  (j2R  ]r�T  (h	h�e]r�T  (hh�eeee]r�T  (hheee]r�T  (jYF  ]r�T  (j[F  ]r�T  (j]F  ]r�T  (h	j�  e]r�T  (hh�e]r�T  (hhe]r�T  (jdF  ]r�T  (h	he]r�T  (hh�e]r�T  (hhe]r�T  (j2R  ]r�T  (h	h�e]r�T  (hh�eeee]r�T  (hheeej�T  j�T  ]r�T  (jYF  ]r�T  (j[F  ]r�T  (j]F  ]r�T  (h	j�  e]r�T  (hh�e]r�T  (hhe]r�T  (jdF  ]r�T  (h	he]r�T  (hh�e]r�T  (hhe]r�T  (j2R  ]r�T  (h	h�e]r�T  (hh�eeee]r�T  (hheeej�T  j�T  j�T  j�T  j�T  j�T  j�T  j�T  j�T  j�T  j�T  j�T  j�T  j�T  j�T  ]r�T  (jYF  ]r�T  (j[F  ]r�T  (j]F  ]r�T  (h	j�  e]r�T  (hh�e]r�T  (hhe]r�T  (jdF  ]r�T  (h	he]r�T  (hh�e]r�T  (hhe]r�T  (j2R  ]r�T  (h	h�e]r�T  (hh�eeee]r�T  (hheeej�T  j�T  j�T  ]r�T  (jYF  ]r�T  (j[F  ]r�T  (j]F  ]r�T  (h	j�  e]r�T  (hh�e]r�T  (hhe]r�T  (jdF  ]r�T  (h	he]r�T  (hh�e]r�T  (hhe]r�T  (j2R  ]r�T  (h	h�e]r�T  (hh�eeee]r�T  (hheeej�T  j�T  j�T  j�T  j�T  ]r U  (jYF  ]rU  (j[F  ]rU  (j]F  ]rU  (h	j�  e]rU  (hh�e]rU  (hhe]rU  (jdF  ]rU  (h	he]rU  (hh�e]r	U  (hhe]r
U  (j2R  ]rU  (h	h�e]rU  (hh�eeee]rU  (hheeej U  j U  j U  j U  j U  ]rU  (jYF  ]rU  (j[F  ]rU  (j]F  ]rU  (h	j�  e]rU  (hh�e]rU  (hhe]rU  (jdF  ]rU  (h	he]rU  (hh�e]rU  (hhe]rU  (j2R  ]rU  (h	h�e]rU  (hh�eeee]rU  (hheeejU  jU  jU  jU  jU  jU  ]rU  (jYF  ]rU  (j[F  ]rU  (j]F  ]rU  (h	j�  e]r U  (hh�e]r!U  (hhe]r"U  (jdF  ]r#U  (h	he]r$U  (hh�e]r%U  (hhe]r&U  (j2R  ]r'U  (h	h�e]r(U  (hh�eeee]r)U  (hheeejU  jU  ]r*U  (jYF  ]r+U  (j[F  ]r,U  (j]F  ]r-U  (h	j�  e]r.U  (hh�e]r/U  (hhe]r0U  (jdF  ]r1U  (h	he]r2U  (hh�e]r3U  (hhe]r4U  (j2R  ]r5U  (h	h�e]r6U  (hh�eeee]r7U  (hheee]r8U  (jYF  ]r9U  (j[F  ]r:U  (j]F  ]r;U  (h	j�  e]r<U  (hh�e]r=U  (hhe]r>U  (jdF  ]r?U  (h	he]r@U  (hh�e]rAU  (hhe]rBU  (j2R  ]rCU  (h	h�e]rDU  (hh�eeee]rEU  (hheeej8U  j8U  j8U  ]rFU  (jYF  ]rGU  (j[F  ]rHU  (j]F  ]rIU  (h	j�  e]rJU  (hh�e]rKU  (hhe]rLU  (jdF  ]rMU  (h	he]rNU  (hh�e]rOU  (hhe]rPU  (j2R  ]rQU  (h	h�e]rRU  (hh�eeee]rSU  (hheeejFU  jFU  jFU  ]rTU  (jYF  ]rUU  (j[F  ]rVU  (j]F  ]rWU  (h	j�  e]rXU  (hh�e]rYU  (hhe]rZU  (jdF  ]r[U  (h	he]r\U  (hh�e]r]U  (hhe]r^U  (j2R  ]r_U  (h	h�e]r`U  (hh�eeee]raU  (hheeejTU  jTU  ]rbU  (jYF  ]rcU  (j[F  ]rdU  (j]F  ]reU  (h	j�  e]rfU  (hh�e]rgU  (hhe]rhU  (jdF  ]riU  (h	he]rjU  (hh�e]rkU  (hhe]rlU  (j2R  ]rmU  (h	h�e]rnU  (hh�eeee]roU  (hheeejbU  jbU  ]rpU  (jYF  ]rqU  (j[F  ]rrU  (j]F  ]rsU  (h	j�  e]rtU  (hh�e]ruU  (hhe]rvU  (jdF  ]rwU  (h	he]rxU  (hh�e]ryU  (hhe]rzU  (j2R  ]r{U  (h	h�e]r|U  (hh�eeee]r}U  (hheeejpU  jpU  ]r~U  (jYF  ]rU  (j[F  ]r�U  (j]F  ]r�U  (h	j�  e]r�U  (hh�e]r�U  (hhe]r�U  (jdF  ]r�U  (h	he]r�U  (hh�e]r�U  (hhe]r�U  (j2R  ]r�U  (h	h�e]r�U  (hh�eeee]r�U  (hheeej~U  j~U  j~U  j~U  j~U  j~U  j~U  ]r�U  (jYF  ]r�U  (j[F  ]r�U  (j]F  ]r�U  (h	j�  e]r�U  (hh�e]r�U  (hhe]r�U  (jdF  ]r�U  (h	he]r�U  (hh�e]r�U  (hhe]r�U  (j2R  ]r�U  (h	h�e]r�U  (hh�eeee]r�U  (hheee]r�U  (jYF  ]r�U  (j[F  ]r�U  (j]F  ]r�U  (h	j�  e]r�U  (hh�e]r�U  (hhe]r�U  (jdF  ]r�U  (h	he]r�U  (hh�e]r�U  (hhe]r�U  (j2R  ]r�U  (h	h�e]r�U  (hh�eeee]r�U  (hheeej�U  j�U  j�U  ]r�U  (jYF  ]r�U  (j[F  ]r�U  (j]F  ]r�U  (h	j�  e]r�U  (hh�e]r�U  (hhe]r�U  (jdF  ]r�U  (h	he]r�U  (hh�e]r�U  (hhe]r�U  (j2R  ]r�U  (h	h�e]r�U  (hh�eeee]r�U  (hheeej�U  ]r�U  (jYF  ]r�U  (j[F  ]r�U  (j]F  ]r�U  (h	j�  e]r�U  (hh�e]r�U  (hhe]r�U  (jdF  ]r�U  (h	he]r�U  (hh�e]r�U  (hhe]r�U  (j2R  ]r�U  (h	h�e]r�U  (hh�eeee]r�U  (hheeej�U  j�U  j�U  j�U  j�U  ]r�U  (jYF  ]r�U  (j[F  ]r�U  (j]F  ]r�U  (h	j�  e]r�U  (hh�e]r�U  (hhe]r�U  (jdF  ]r�U  (h	he]r�U  (hh�e]r�U  (hhe]r�U  (j2R  ]r�U  (h	h�e]r�U  (hh�eeee]r�U  (hheee]r�U  (jYF  ]r�U  (j[F  ]r�U  (j]F  ]r�U  (h	j�  e]r�U  (hh�e]r�U  (hhe]r�U  (jdF  ]r�U  (h	he]r�U  (hh�e]r�U  (hhe]r�U  (j2R  ]r�U  (h	h�e]r�U  (hh�eeee]r�U  (hheeej�U  j�U  j�U  j�U  j�U  j�U  j�U  j�U  ]r�U  (jYF  ]r�U  (j[F  ]r�U  (j]F  ]r�U  (h	j�  e]r�U  (hh�e]r�U  (hhe]r�U  (jdF  ]r�U  (h	he]r�U  (hh�e]r�U  (hhe]r�U  (j2R  ]r�U  (h	h�e]r�U  (hh�eeee]r�U  (hheeej�U  j�U  j�U  j�U  j�U  ]r�U  (jYF  ]r�U  (j[F  ]r�U  (j]F  ]r�U  (h	j�  e]r�U  (hh�e]r�U  (hhe]r�U  (jdF  ]r�U  (h	he]r�U  (hh�e]r�U  (hhe]r�U  (j2R  ]r�U  (h	h�e]r�U  (hh�eeee]r�U  (hheeej�U  j�U  j�U  j�U  ]r�U  (jYF  ]r�U  (j[F  ]r�U  (j]F  ]r�U  (h	j�  e]r V  (hh�e]rV  (hhe]rV  (jdF  ]rV  (h	he]rV  (hh�e]rV  (hhe]rV  (j2R  ]rV  (h	h�e]rV  (hh�eeee]r	V  (hheee]r
V  (jYF  ]rV  (j[F  ]rV  (j]F  ]rV  (h	j�  e]rV  (hh�e]rV  (hhe]rV  (jdF  ]rV  (h	he]rV  (hh�e]rV  (hhe]rV  (j2R  ]rV  (h	h�e]rV  (hh�eeee]rV  (hheee]rV  (jYF  ]rV  (j[F  ]rV  (j]F  ]rV  (h	j�  e]rV  (hh�e]rV  (hhe]rV  (jdF  ]rV  (h	he]r V  (hh�e]r!V  (hhe]r"V  (j2R  ]r#V  (h	h�e]r$V  (hh�eeee]r%V  (hheeejV  ]r&V  (jYF  ]r'V  (j[F  ]r(V  (j]F  ]r)V  (h	j�  e]r*V  (hh�e]r+V  (hhe]r,V  (jdF  ]r-V  (h	he]r.V  (hh�e]r/V  (hhe]r0V  (j2R  ]r1V  (h	h�e]r2V  (hh�eeee]r3V  (hheeej&V  j&V  j&V  j&V  j&V  ]r4V  (jYF  ]r5V  (j[F  ]r6V  (j]F  ]r7V  (h	j�  e]r8V  (hh�e]r9V  (hhe]r:V  (jdF  ]r;V  (h	he]r<V  (hh�e]r=V  (hhe]r>V  (j2R  ]r?V  (h	h�e]r@V  (hh�eeee]rAV  (hheee]rBV  (jYF  ]rCV  (j[F  ]rDV  (j]F  ]rEV  (h	j�  e]rFV  (hh�e]rGV  (hhe]rHV  (jdF  ]rIV  (h	he]rJV  (hh�e]rKV  (hhe]rLV  (j2R  ]rMV  (h	h�e]rNV  (hh�eeee]rOV  (hheee]rPV  (jYF  ]rQV  (j[F  ]rRV  (j]F  ]rSV  (h	j�  e]rTV  (hh�e]rUV  (hhe]rVV  (jdF  ]rWV  (h	he]rXV  (hh�e]rYV  (hhe]rZV  (j2R  ]r[V  (h	h�e]r\V  (hh�eeee]r]V  (hheeejPV  jPV  jPV  ]r^V  (jYF  ]r_V  (j[F  ]r`V  (j]F  ]raV  (h	j�  e]rbV  (hh�e]rcV  (hhe]rdV  (jdF  ]reV  (h	he]rfV  (hh�e]rgV  (hhe]rhV  (j2R  ]riV  (h	h�e]rjV  (hh�eeee]rkV  (hheeej^V  ]rlV  (jYF  ]rmV  (j[F  ]rnV  (j]F  ]roV  (h	j�  e]rpV  (hh�e]rqV  (hhe]rrV  (jdF  ]rsV  (h	he]rtV  (hh�e]ruV  (hhe]rvV  (j2R  ]rwV  (h	h�e]rxV  (hh�eeee]ryV  (hheeejlV  ]rzV  (jYF  ]r{V  (j[F  ]r|V  (j]F  ]r}V  (h	j�  e]r~V  (hh�e]rV  (hhe]r�V  (jdF  ]r�V  (h	he]r�V  (hh�e]r�V  (hhe]r�V  (j2R  ]r�V  (h	h�e]r�V  (hh�eeee]r�V  (hheeejzV  jzV  jzV  jzV  ]r�V  (jYF  ]r�V  (j[F  ]r�V  (j]F  ]r�V  (h	j�  e]r�V  (hh�e]r�V  (hhe]r�V  (jdF  ]r�V  (h	he]r�V  (hh�e]r�V  (hhe]r�V  (j2R  ]r�V  (h	h�e]r�V  (hh�eeee]r�V  (hheeej�V  j�V  ]r�V  (jYF  ]r�V  (j[F  ]r�V  (j]F  ]r�V  (h	j�  e]r�V  (hh�e]r�V  (hhe]r�V  (jdF  ]r�V  (h	he]r�V  (hh�e]r�V  (hhe]r�V  (j2R  ]r�V  (h	h�e]r�V  (hh�eeee]r�V  (hheeej�V  j�V  ]r�V  (jYF  ]r�V  (j[F  ]r�V  (j]F  ]r�V  (h	j�  e]r�V  (hh�e]r�V  (hhe]r�V  (jdF  ]r�V  (h	he]r�V  (hh�e]r�V  (hhe]r�V  (j2R  ]r�V  (h	h�e]r�V  (hh�eeee]r�V  (hheeej�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  ]r�V  (jYF  ]r�V  (j[F  ]r�V  (j]F  ]r�V  (h	j�  e]r�V  (hh�e]r�V  (hhe]r�V  (jdF  ]r�V  (h	he]r�V  (hh�e]r�V  (hhe]r�V  (j2R  ]r�V  (h	h�e]r�V  (hh�eeee]r�V  (hheee]r�V  (jYF  ]r�V  (j[F  ]r�V  (j]F  ]r�V  (h	j�  e]r�V  (hh�e]r�V  (hhe]r�V  (jdF  ]r�V  (h	he]r�V  (hh�e]r�V  (hhe]r�V  (j2R  ]r�V  (h	h�e]r�V  (hh�eeee]r�V  (hheeej�V  j�V  j�V  ]r�V  (jYF  ]r�V  (j[F  ]r�V  (j]F  ]r�V  (h	j�  e]r�V  (hh�e]r�V  (hhe]r�V  (jdF  ]r�V  (h	he]r�V  (hh�e]r�V  (hhe]r�V  (j2R  ]r�V  (h	h�e]r�V  (hh�eeee]r�V  (hheeej�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  ]r�V  (jYF  ]r�V  (j[F  ]r�V  (j]F  ]r�V  (h	j�  e]r�V  (hh�e]r�V  (hhe]r�V  (jdF  ]r�V  (h	he]r�V  (hh�e]r�V  (hhe]r�V  (j2R  ]r�V  (h	h�e]r�V  (hh�eeee]r�V  (hheeej�V  j�V  ]r�V  (jYF  ]r�V  (j[F  ]r�V  (j]F  ]r�V  (h	j�  e]r�V  (hh�e]r�V  (hhe]r�V  (jdF  ]r�V  (h	he]r�V  (hh�e]r�V  (hhe]r�V  (j2R  ]r�V  (h	h�e]r�V  (hh�eeee]r�V  (hheeej�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  j�V  ]r�V  (jYF  ]r�V  (j[F  ]r�V  (j]F  ]r�V  (h	j�  e]r�V  (hh�e]r�V  (hhe]r�V  (jdF  ]r�V  (h	he]r W  (hh�e]rW  (hhe]rW  (j2R  ]rW  (h	h�e]rW  (hh�eeee]rW  (hheee]rW  (jYF  ]rW  (j[F  ]rW  (j]F  ]r	W  (h	j�  e]r
W  (hh�e]rW  (hhe]rW  (jdF  ]rW  (h	he]rW  (hh�e]rW  (hhe]rW  (j2R  ]rW  (h	h�e]rW  (hh�eeee]rW  (hheeejW  jW  jW  ]rW  (jYF  ]rW  (j[F  ]rW  (j]F  ]rW  (h	j�  e]rW  (hh�e]rW  (hhe]rW  (jdF  ]rW  (h	he]rW  (hh�e]rW  (hhe]rW  (j2R  ]rW  (h	h�e]r W  (hh�eeee]r!W  (hheeejW  jW  jW  jW  jW  jW  ]r"W  (jYF  ]r#W  (j[F  ]r$W  (j]F  ]r%W  (h	j�  e]r&W  (hh�e]r'W  (hhe]r(W  (jdF  ]r)W  (h	he]r*W  (hh�e]r+W  (hhe]r,W  (j2R  ]r-W  (h	h�e]r.W  (hh�eeee]r/W  (hheeej"W  ]r0W  (jYF  ]r1W  (j[F  ]r2W  (j]F  ]r3W  (h	j�  e]r4W  (hh�e]r5W  (hhe]r6W  (jdF  ]r7W  (h	he]r8W  (hh�e]r9W  (hhe]r:W  (j2R  ]r;W  (h	h�e]r<W  (hh�eeee]r=W  (hheeej0W  j0W  ]r>W  (jYF  ]r?W  (j[F  ]r@W  (j]F  ]rAW  (h	j�  e]rBW  (hh�e]rCW  (hhe]rDW  (jdF  ]rEW  (h	he]rFW  (hh�e]rGW  (hhe]rHW  (j2R  ]rIW  (h	h�e]rJW  (hh�eeee]rKW  (hheeej>W  j>W  j>W  j>W  ]rLW  (jYF  ]rMW  (j[F  ]rNW  (j]F  ]rOW  (h	j�  e]rPW  (hh�e]rQW  (hhe]rRW  (jdF  ]rSW  (h	he]rTW  (hh�e]rUW  (hhe]rVW  (j2R  ]rWW  (h	h�e]rXW  (hh�eeee]rYW  (hheeejLW  ]rZW  (jYF  ]r[W  (j[F  ]r\W  (j]F  ]r]W  (h	j�  e]r^W  (hh�e]r_W  (hhe]r`W  (jdF  ]raW  (h	he]rbW  (hh�e]rcW  (hhe]rdW  (j2R  ]reW  (h	h�e]rfW  (hh�eeee]rgW  (hheeejZW  jZW  jZW  jZW  jZW  jZW  jZW  jZW  jZW  jZW  jZW  jZW  ]rhW  (jYF  ]riW  (j[F  ]rjW  (j]F  ]rkW  (h	j�  e]rlW  (hh�e]rmW  (hhe]rnW  (jdF  ]roW  (h	he]rpW  (hh�e]rqW  (hhe]rrW  (j2R  ]rsW  (h	h�e]rtW  (hh�eeee]ruW  (hheee]rvW  (jYF  ]rwW  (j[F  ]rxW  (j]F  ]ryW  (h	j�  e]rzW  (hh�e]r{W  (hhe]r|W  (jdF  ]r}W  (h	he]r~W  (hh�e]rW  (hhe]r�W  (j2R  ]r�W  (h	h�e]r�W  (hh�eeee]r�W  (hheeejvW  jvW  jvW  jvW  jvW  jvW  jvW  ]r�W  (jYF  ]r�W  (j[F  ]r�W  (j]F  ]r�W  (h	j�  e]r�W  (hh�e]r�W  (hhe]r�W  (jdF  ]r�W  (h	he]r�W  (hh�e]r�W  (hhe]r�W  (j2R  ]r�W  (h	h�e]r�W  (hh�eeee]r�W  (hheee]r�W  (jYF  ]r�W  (j[F  ]r�W  (j]F  ]r�W  (h	j�  e]r�W  (hh�e]r�W  (hhe]r�W  (jdF  ]r�W  (h	he]r�W  (hh�e]r�W  (hhe]r�W  (j2R  ]r�W  (h	h�e]r�W  (hh�eeee]r�W  (hheeej�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  ]r�W  (jYF  ]r�W  (j[F  ]r�W  (j]F  ]r�W  (h	j�  e]r�W  (hh�e]r�W  (hhe]r�W  (jdF  ]r�W  (h	he]r�W  (hh�e]r�W  (hhe]r�W  (j2R  ]r�W  (h	h�e]r�W  (hh�eeee]r�W  (hheeej�W  ]r�W  (jYF  ]r�W  (j[F  ]r�W  (j]F  ]r�W  (h	j�  e]r�W  (hh�e]r�W  (hhe]r�W  (jdF  ]r�W  (h	he]r�W  (hh�e]r�W  (hhe]r�W  (j2R  ]r�W  (h	h�e]r�W  (hh�eeee]r�W  (hheeej�W  j�W  j�W  j�W  j�W  j�W  ]r�W  (jYF  ]r�W  (j[F  ]r�W  (j]F  ]r�W  (h	j�  e]r�W  (hh�e]r�W  (hhe]r�W  (jdF  ]r�W  (h	he]r�W  (hh�e]r�W  (hhe]r�W  (j2R  ]r�W  (h	h�e]r�W  (hh�eeee]r�W  (hheeej�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  j�W  ]r�W  (jYF  ]r�W  (j[F  ]r�W  (j]F  ]r�W  (h	j�  e]r�W  (hh�e]r�W  (hhe]r�W  (jdF  ]r�W  (h	he]r�W  (hh�e]r�W  (hhe]r�W  (j2R  ]r�W  (h	h�e]r�W  (hh�eeee]r�W  (hheee]r�W  (jYF  ]r�W  (j[F  ]r�W  (j]F  ]r�W  (h	j�  e]r�W  (hh�e]r�W  (hhe]r�W  (jdF  ]r�W  (h	he]r�W  (hh�e]r�W  (hhe]r�W  (j2R  ]r�W  (h	h�e]r�W  (hh�eeee]r�W  (hheee]r�W  (jYF  ]r�W  (j[F  ]r�W  (j]F  ]r�W  (h	j�  e]r�W  (hh�e]r�W  (hhe]r�W  (jdF  ]r�W  (h	he]r�W  (hh�e]r�W  (hhe]r�W  (j2R  ]r�W  (h	h�e]r�W  (hh�eeee]r�W  (hheeej�W  j�W  ]r�W  (jYF  ]r�W  (j[F  ]r�W  (j]F  ]r�W  (h	j�  e]r�W  (hh�e]r�W  (hhe]r�W  (jdF  ]r�W  (h	he]r�W  (hh�e]r�W  (hhe]r�W  (j2R  ]r�W  (h	h�e]r X  (hh�eeee]rX  (hheeej�W  j�W  j�W  ]rX  (jYF  ]rX  (j[F  ]rX  (j]F  ]rX  (h	j�  e]rX  (hh�e]rX  (hhe]rX  (jdF  ]r	X  (h	he]r
X  (hh�e]rX  (hhe]rX  (j2R  ]rX  (h	h�e]rX  (hh�eeee]rX  (hheeejX  jX  ]rX  (jYF  ]rX  (j[F  ]rX  (j]F  ]rX  (h	j�  e]rX  (hh�e]rX  (hhe]rX  (jdF  ]rX  (h	he]rX  (hh�e]rX  (hhe]rX  (j2R  ]rX  (h	h�e]rX  (hh�eeee]rX  (hheeejX  jX  jX  jX  jX  jX  jX  ]rX  (jYF  ]rX  (j[F  ]r X  (j]F  ]r!X  (h	j�  e]r"X  (hh�e]r#X  (hhe]r$X  (jdF  ]r%X  (h	he]r&X  (hh�e]r'X  (hhe]r(X  (j2R  ]r)X  (h	h�e]r*X  (hh�eeee]r+X  (hheeejX  jX  jX  jX  jX  jX  jX  jX  jX  jX  ]r,X  (jYF  ]r-X  (j[F  ]r.X  (j]F  ]r/X  (h	j�  e]r0X  (hh�e]r1X  (hhe]r2X  (jdF  ]r3X  (h	he]r4X  (hh�e]r5X  (hhe]r6X  (j2R  ]r7X  (h	h�e]r8X  (hh�eeee]r9X  (hheeej,X  j,X  j,X  j,X  j,X  ]r:X  (jYF  ]r;X  (j[F  ]r<X  (j]F  ]r=X  (h	j�  e]r>X  (hh�e]r?X  (hhe]r@X  (jdF  ]rAX  (h	he]rBX  (hh�e]rCX  (hhe]rDX  (j2R  ]rEX  (h	h�e]rFX  (hh�eeee]rGX  (hheeej:X  j:X  j:X  j:X  j:X  j:X  j:X  j:X  j:X  j:X  j:X  j:X  ]rHX  (jYF  ]rIX  (j[F  ]rJX  (j]F  ]rKX  (h	j�  e]rLX  (hh�e]rMX  (hhe]rNX  (jdF  ]rOX  (h	he]rPX  (hh�e]rQX  (hhe]rRX  (j2R  ]rSX  (h	h�e]rTX  (hh�eeee]rUX  (hheeejHX  jHX  jHX  jHX  jHX  jHX  jHX  jHX  ]rVX  (jYF  ]rWX  (j[F  ]rXX  (j]F  ]rYX  (h	j�  e]rZX  (hh�e]r[X  (hhe]r\X  (jdF  ]r]X  (h	he]r^X  (hh�e]r_X  (hhe]r`X  (j2R  ]raX  (h	h�e]rbX  (hh�eeee]rcX  (hheeejVX  jVX  ]rdX  (jYF  ]reX  (j[F  ]rfX  (j]F  ]rgX  (h	j�  e]rhX  (hh�e]riX  (hhe]rjX  (jdF  ]rkX  (h	he]rlX  (hh�e]rmX  (hhe]rnX  (j2R  ]roX  (h	h�e]rpX  (hh�eeee]rqX  (hheeejdX  jdX  jdX  ]rrX  (jYF  ]rsX  (j[F  ]rtX  (j]F  ]ruX  (h	j�  e]rvX  (hh�e]rwX  (hhe]rxX  (jdF  ]ryX  (h	he]rzX  (hh�e]r{X  (hhe]r|X  (j2R  ]r}X  (h	h�e]r~X  (hh�eeee]rX  (hheeejrX  ]r�X  (jYF  ]r�X  (j[F  ]r�X  (j]F  ]r�X  (h	j�  e]r�X  (hh�e]r�X  (hhe]r�X  (jdF  ]r�X  (h	he]r�X  (hh�e]r�X  (hhe]r�X  (j2R  ]r�X  (h	h�e]r�X  (hh�eeee]r�X  (hheeej�X  ]r�X  (jYF  ]r�X  (j[F  ]r�X  (j]F  ]r�X  (h	j�  e]r�X  (hh�e]r�X  (hhe]r�X  (jdF  ]r�X  (h	he]r�X  (hh�e]r�X  (hhe]r�X  (j2R  ]r�X  (h	h�e]r�X  (hh�eeee]r�X  (hheeej�X  j�X  j�X  ]r�X  (jYF  ]r�X  (j[F  ]r�X  (j]F  ]r�X  (h	j�  e]r�X  (hh�e]r�X  (hhe]r�X  (jdF  ]r�X  (h	he]r�X  (hh�e]r�X  (hhe]r�X  (j2R  ]r�X  (h	h�e]r�X  (hh�eeee]r�X  (hheee]r�X  (jYF  ]r�X  (j[F  ]r�X  (j]F  ]r�X  (h	j�  e]r�X  (hh�e]r�X  (hhe]r�X  (jdF  ]r�X  (h	he]r�X  (hh�e]r�X  (hhe]r�X  (j2R  ]r�X  (h	h�e]r�X  (hh�eeee]r�X  (hheeej�X  j�X  j�X  j�X  j�X  j�X  ]r�X  (jYF  ]r�X  (j[F  ]r�X  (j]F  ]r�X  (h	j�  e]r�X  (hh�e]r�X  (hhe]r�X  (jdF  ]r�X  (h	he]r�X  (hh�e]r�X  (hhe]r�X  (j2R  ]r�X  (h	h�e]r�X  (hh�eeee]r�X  (hheeej�X  j�X  j�X  j�X  ]r�X  (jYF  ]r�X  (j[F  ]r�X  (j]F  ]r�X  (h	j�  e]r�X  (hh�e]r�X  (hhe]r�X  (jdF  ]r�X  (h	he]r�X  (hh�e]r�X  (hhe]r�X  (j2R  ]r�X  (h	h�e]r�X  (hh�eeee]r�X  (hheee]r�X  (jYF  ]r�X  (j[F  ]r�X  (j]F  ]r�X  (h	j�  e]r�X  (hh�e]r�X  (hhe]r�X  (jdF  ]r�X  (h	he]r�X  (hh�e]r�X  (hhe]r�X  (j2R  ]r�X  (h	h�e]r�X  (hh�eeee]r�X  (hheeej�X  j�X  ]r�X  (jYF  ]r�X  (j[F  ]r�X  (j]F  ]r�X  (h	j�  e]r�X  (hh�e]r�X  (hhe]r�X  (jdF  ]r�X  (h	he]r�X  (hh�e]r�X  (hhe]r�X  (j2R  ]r�X  (h	h�e]r�X  (hh�eeee]r�X  (hheeej�X  ]r�X  (jYF  ]r�X  (j[F  ]r�X  (j]F  ]r�X  (h	j�  e]r�X  (hh�e]r�X  (hhe]r�X  (jdF  ]r�X  (h	he]r�X  (hh�e]r�X  (hhe]r�X  (j2R  ]r�X  (h	h�e]r�X  (hh�eeee]r�X  (hheeej�X  j�X  j�X  j�X  j�X  j�X  j�X  j�X  ]r�X  (jYF  ]r�X  (j[F  ]r Y  (j]F  ]rY  (h	j�  e]rY  (hh�e]rY  (hhe]rY  (jdF  ]rY  (h	he]rY  (hh�e]rY  (hhe]rY  (j2R  ]r	Y  (h	h�e]r
Y  (hh�eeee]rY  (hheeej�X  j�X  j�X  ]rY  (jYF  ]rY  (j[F  ]rY  (j]F  ]rY  (h	j�  e]rY  (hh�e]rY  (hhe]rY  (jdF  ]rY  (h	he]rY  (hh�e]rY  (hhe]rY  (j2R  ]rY  (h	h�e]rY  (hh�eeee]rY  (hheeejY  jY  jY  jY  jY  jY  ]rY  (jYF  ]rY  (j[F  ]rY  (j]F  ]rY  (h	j�  e]rY  (hh�e]rY  (hhe]r Y  (jdF  ]r!Y  (h	he]r"Y  (hh�e]r#Y  (hhe]r$Y  (j2R  ]r%Y  (h	h�e]r&Y  (hh�eeee]r'Y  (hheeejY  ]r(Y  (jYF  ]r)Y  (j[F  ]r*Y  (j]F  ]r+Y  (h	j�  e]r,Y  (hh�e]r-Y  (hhe]r.Y  (jdF  ]r/Y  (h	he]r0Y  (hh�e]r1Y  (hhe]r2Y  (j2R  ]r3Y  (h	h�e]r4Y  (hh�eeee]r5Y  (hheeej(Y  j(Y  j(Y  ]r6Y  (jYF  ]r7Y  (j[F  ]r8Y  (j]F  ]r9Y  (h	j�  e]r:Y  (hh�e]r;Y  (hhe]r<Y  (jdF  ]r=Y  (h	he]r>Y  (hh�e]r?Y  (hhe]r@Y  (j2R  ]rAY  (h	h�e]rBY  (hh�eeee]rCY  (hheee]rDY  (jYF  ]rEY  (j[F  ]rFY  (j]F  ]rGY  (h	j�  e]rHY  (hh�e]rIY  (hhe]rJY  (jdF  ]rKY  (h	he]rLY  (hh�e]rMY  (hhe]rNY  (j2R  ]rOY  (h	h�e]rPY  (hh�eeee]rQY  (hheeejDY  jDY  jDY  jDY  jDY  jDY  jDY  ]rRY  (jYF  ]rSY  (j[F  ]rTY  (j]F  ]rUY  (h	j�  e]rVY  (hh�e]rWY  (hhe]rXY  (jdF  ]rYY  (h	he]rZY  (hh�e]r[Y  (hhe]r\Y  (j2R  ]r]Y  (h	h�e]r^Y  (hh�eeee]r_Y  (hheee]r`Y  (jYF  ]raY  (j[F  ]rbY  (j]F  ]rcY  (h	j�  e]rdY  (hh�e]reY  (hhe]rfY  (jdF  ]rgY  (h	he]rhY  (hh�e]riY  (hhe]rjY  (j2R  ]rkY  (h	h�e]rlY  (hh�eeee]rmY  (hheee]rnY  (jYF  ]roY  (j[F  ]rpY  (j]F  ]rqY  (h	j�  e]rrY  (hh�e]rsY  (hhe]rtY  (jdF  ]ruY  (h	he]rvY  (hh�e]rwY  (hhe]rxY  (j2R  ]ryY  (h	h�e]rzY  (hh�eeee]r{Y  (hheee]r|Y  (jYF  ]r}Y  (j[F  ]r~Y  (j]F  ]rY  (h	j�  e]r�Y  (hh�e]r�Y  (hhe]r�Y  (jdF  ]r�Y  (h	he]r�Y  (hh�e]r�Y  (hhe]r�Y  (j2R  ]r�Y  (h	h�e]r�Y  (hh�eeee]r�Y  (hheeej|Y  j|Y  ]r�Y  (jYF  ]r�Y  (j[F  ]r�Y  (j]F  ]r�Y  (h	j�  e]r�Y  (hh�e]r�Y  (hhe]r�Y  (jdF  ]r�Y  (h	he]r�Y  (hh�e]r�Y  (hhe]r�Y  (j2R  ]r�Y  (h	h�e]r�Y  (hh�eeee]r�Y  (hheeej�Y  ]r�Y  (jYF  ]r�Y  (j[F  ]r�Y  (j]F  ]r�Y  (h	j�  e]r�Y  (hh�e]r�Y  (hhe]r�Y  (jdF  ]r�Y  (h	he]r�Y  (hh�e]r�Y  (hhe]r�Y  (j2R  ]r�Y  (h	h�e]r�Y  (hh�eeee]r�Y  (hheeej�Y  j�Y  j�Y  j�Y  j�Y  j�Y  j�Y  ]r�Y  (jYF  ]r�Y  (j[F  ]r�Y  (j]F  ]r�Y  (h	j�  e]r�Y  (hh�e]r�Y  (hhe]r�Y  (jdF  ]r�Y  (h	he]r�Y  (hh�e]r�Y  (hhe]r�Y  (j2R  ]r�Y  (h	h�e]r�Y  (hh�eeee]r�Y  (hheee]r�Y  (jYF  ]r�Y  (j[F  ]r�Y  (j]F  ]r�Y  (h	h�e]r�Y  (hh�e]r�Y  (hhe]r�Y  (jdF  ]r�Y  (h	he]r�Y  (hh�e]r�Y  (hhe]r�Y  (j2R  ]r�Y  (h	h�e]r�Y  (hh�eeee]r�Y  (hheeej�Y  j�Y  ]r�Y  (jYF  ]r�Y  (j[F  ]r�Y  (j]F  ]r�Y  (h	h�e]r�Y  (hh�e]r�Y  (hhe]r�Y  (jdF  ]r�Y  (h	he]r�Y  (hh�e]r�Y  (hhe]r�Y  (j2R  ]r�Y  (h	h�e]r�Y  (hh�eeee]r�Y  (hheeej�Y  ]r�Y  (jYF  ]r�Y  (j[F  ]r�Y  (j]F  ]r�Y  (h	h�e]r�Y  (hh�e]r�Y  (hhe]r�Y  (jdF  ]r�Y  (h	he]r�Y  (hh�e]r�Y  (hhe]r�Y  (j2R  ]r�Y  (h	h�e]r�Y  (hh�eeee]r�Y  (hheeej�Y  ]r�Y  (jYF  ]r�Y  (j[F  ]r�Y  (j]F  ]r�Y  (h	h�e]r�Y  (hh�e]r�Y  (hhe]r�Y  (jdF  ]r�Y  (h	he]r�Y  (hh�e]r�Y  (hhe]r�Y  (j2R  ]r�Y  (h	h�e]r�Y  (hh�eeee]r�Y  (hheeej�Y  j�Y  j�Y  j�Y  j�Y  j�Y  ]r�Y  (jYF  ]r�Y  (j[F  ]r�Y  (j]F  ]r�Y  (h	h�e]r�Y  (hh�e]r�Y  (hhe]r�Y  (jdF  ]r�Y  (h	he]r�Y  (hh�e]r�Y  (hhe]r�Y  (j2R  ]r�Y  (h	h�e]r�Y  (hh�eeee]r�Y  (hheeej�Y  j�Y  ]r�Y  (jYF  ]r�Y  (j[F  ]r�Y  (j]F  ]r�Y  (h	h�e]r�Y  (hh�e]r�Y  (hhe]r Z  (jdF  ]rZ  (h	he]rZ  (hh�e]rZ  (hhe]rZ  (j2R  ]rZ  (h	h�e]rZ  (hh�eeee]rZ  (hheeej�Y  j�Y  j�Y  j�Y  j�Y  j�Y  j�Y  j�Y  j�Y  j�Y  j�Y  j�Y  j�Y  ]rZ  (jYF  ]r	Z  (j[F  ]r
Z  (j]F  ]rZ  (h	j�  e]rZ  (hh�e]rZ  (hhe]rZ  (jdF  ]rZ  (h	he]rZ  (hh�e]rZ  (hhe]rZ  (j2R  ]rZ  (h	h�e]rZ  (hh�eeee]rZ  (hheeejZ  jZ  jZ  jZ  jZ  ]rZ  (jYF  ]rZ  (j[F  ]rZ  (j]F  ]rZ  (h	j�  e]rZ  (hh�e]rZ  (hhe]rZ  (jdF  ]rZ  (h	he]rZ  (hh�e]rZ  (hhe]r Z  (j2R  ]r!Z  (h	h�e]r"Z  (hh�eeee]r#Z  (hheee]r$Z  (jYF  ]r%Z  (j[F  ]r&Z  (j]F  ]r'Z  (h	j�  e]r(Z  (hh�e]r)Z  (hhe]r*Z  (jdF  ]r+Z  (h	he]r,Z  (hh�e]r-Z  (hhe]r.Z  (j2R  ]r/Z  (h	h�e]r0Z  (hh�eeee]r1Z  (hheeej$Z  ]r2Z  (jYF  ]r3Z  (j[F  ]r4Z  (j]F  ]r5Z  (h	j�  e]r6Z  (hh�e]r7Z  (hhe]r8Z  (jdF  ]r9Z  (h	he]r:Z  (hh�e]r;Z  (hhe]r<Z  (j2R  ]r=Z  (h	h�e]r>Z  (hh�eeee]r?Z  (hheeej2Z  j2Z  j2Z  j2Z  j2Z  j2Z  ]r@Z  (jYF  ]rAZ  (j[F  ]rBZ  (j]F  ]rCZ  (h	j�  e]rDZ  (hh�e]rEZ  (hhe]rFZ  (jdF  ]rGZ  (h	he]rHZ  (hh�e]rIZ  (hhe]rJZ  (j2R  ]rKZ  (h	h�e]rLZ  (hh�eeee]rMZ  (hheeej@Z  j@Z  j@Z  j@Z  ]rNZ  (jYF  ]rOZ  (j[F  ]rPZ  (j]F  ]rQZ  (h	j�  e]rRZ  (hh�e]rSZ  (hhe]rTZ  (jdF  ]rUZ  (h	he]rVZ  (hh�e]rWZ  (hhe]rXZ  (j2R  ]rYZ  (h	h�e]rZZ  (hh�eeee]r[Z  (hheee]r\Z  (jYF  ]r]Z  (j[F  ]r^Z  (j]F  ]r_Z  (h	j�  e]r`Z  (hh�e]raZ  (hhe]rbZ  (jdF  ]rcZ  (h	he]rdZ  (hh�e]reZ  (hhe]rfZ  (j2R  ]rgZ  (h	h�e]rhZ  (hh�eeee]riZ  (hheee]rjZ  (jYF  ]rkZ  (j[F  ]rlZ  (j]F  ]rmZ  (h	j�  e]rnZ  (hh�e]roZ  (hhe]rpZ  (jdF  ]rqZ  (h	he]rrZ  (hh�e]rsZ  (hhe]rtZ  (j2R  ]ruZ  (h	h�e]rvZ  (hh�eeee]rwZ  (hheeejjZ  jjZ  jjZ  jjZ  jjZ  jjZ  jjZ  jjZ  jjZ  jjZ  jjZ  jjZ  ]rxZ  (jYF  ]ryZ  (j[F  ]rzZ  (j]F  ]r{Z  (h	j�  e]r|Z  (hh�e]r}Z  (hhe]r~Z  (jdF  ]rZ  (h	he]r�Z  (hh�e]r�Z  (hhe]r�Z  (j2R  ]r�Z  (h	h�e]r�Z  (hh�eeee]r�Z  (hheeejxZ  jxZ  jxZ  jxZ  ]r�Z  (jYF  ]r�Z  (j[F  ]r�Z  (j]F  ]r�Z  (h	j�  e]r�Z  (hh�e]r�Z  (hhe]r�Z  (jdF  ]r�Z  (h	he]r�Z  (hh�e]r�Z  (hhe]r�Z  (j2R  ]r�Z  (h	h�e]r�Z  (hh�eeee]r�Z  (hheeej�Z  j�Z  ]r�Z  (jYF  ]r�Z  (j[F  ]r�Z  (j]F  ]r�Z  (h	j�  e]r�Z  (hh�e]r�Z  (hhe]r�Z  (jdF  ]r�Z  (h	he]r�Z  (hh�e]r�Z  (hhe]r�Z  (j2R  ]r�Z  (h	h�e]r�Z  (hh�eeee]r�Z  (hheeej�Z  j�Z  j�Z  j�Z  j�Z  j�Z  j�Z  ]r�Z  (jYF  ]r�Z  (j[F  ]r�Z  (j]F  ]r�Z  (h	j�  e]r�Z  (hh�e]r�Z  (hhe]r�Z  (jdF  ]r�Z  (h	he]r�Z  (hh�e]r�Z  (hhe]r�Z  (j2R  ]r�Z  (h	h�e]r�Z  (hh�eeee]r�Z  (hheeej�Z  j�Z  j�Z  ]r�Z  (jYF  ]r�Z  (j[F  ]r�Z  (j]F  ]r�Z  (h	j�  e]r�Z  (hh�e]r�Z  (hhe]r�Z  (jdF  ]r�Z  (h	he]r�Z  (hh�e]r�Z  (hhe]r�Z  (j2R  ]r�Z  (h	h�e]r�Z  (hh�eeee]r�Z  (hheee]r�Z  (jYF  ]r�Z  (j[F  ]r�Z  (j]F  ]r�Z  (h	j�  e]r�Z  (hh�e]r�Z  (hhe]r�Z  (jdF  ]r�Z  (h	he]r�Z  (hh�e]r�Z  (hhe]r�Z  (j2R  ]r�Z  (h	h�e]r�Z  (hh�eeee]r�Z  (hheeej�Z  j�Z  j�Z  ]r�Z  (jYF  ]r�Z  (j[F  ]r�Z  (j]F  ]r�Z  (h	j�  e]r�Z  (hh�e]r�Z  (hhe]r�Z  (jdF  ]r�Z  (h	he]r�Z  (hh�e]r�Z  (hhe]r�Z  (j2R  ]r�Z  (h	h�e]r�Z  (hh�eeee]r�Z  (hheeej�Z  j�Z  j�Z  ]r�Z  (jYF  ]r�Z  (j[F  ]r�Z  (j]F  ]r�Z  (h	j�  e]r�Z  (hh�e]r�Z  (hhe]r�Z  (jdF  ]r�Z  (h	he]r�Z  (hh�e]r�Z  (hhe]r�Z  (j2R  ]r�Z  (h	h�e]r�Z  (hh�eeee]r�Z  (hheeej�Z  j�Z  j�Z  j�Z  j�Z  j�Z  j�Z  j�Z  j�Z  ]r�Z  (jYF  ]r�Z  (j[F  ]r�Z  (j]F  ]r�Z  (h	j�  e]r�Z  (hh�e]r�Z  (hhe]r�Z  (jdF  ]r�Z  (h	he]r�Z  (hh�e]r�Z  (hhe]r�Z  (j2R  ]r�Z  (h	h�e]r�Z  (hh�eeee]r�Z  (hheeej�Z  j�Z  j�Z  ]r�Z  (jYF  ]r�Z  (j[F  ]r�Z  (j]F  ]r�Z  (h	j�  e]r�Z  (hh�e]r�Z  (hhe]r�Z  (jdF  ]r�Z  (h	he]r�Z  (hh�e]r�Z  (hhe]r [  (j2R  ]r[  (h	h�e]r[  (hh�eeee]r[  (hheeej�Z  j�Z  j�Z  j�Z  j�Z  j�Z  ]r[  (jYF  ]r[  (j[F  ]r[  (j]F  ]r[  (h	j�  e]r[  (hh�e]r	[  (hhe]r
[  (jdF  ]r[  (h	he]r[  (hh�e]r[  (hhe]r[  (j2R  ]r[  (h	h�e]r[  (hh�eeee]r[  (hheeej[  j[  ]r[  (jYF  ]r[  (j[F  ]r[  (j]F  ]r[  (h	j�  e]r[  (hh�e]r[  (hhe]r[  (jdF  ]r[  (h	he]r[  (hh�e]r[  (hhe]r[  (j2R  ]r[  (h	h�e]r[  (hh�eeee]r[  (hheeej[  ]r [  (jYF  ]r![  (j[F  ]r"[  (j]F  ]r#[  (h	j�  e]r$[  (hh�e]r%[  (hhe]r&[  (jdF  ]r'[  (h	he]r([  (hh�e]r)[  (hhe]r*[  (j2R  ]r+[  (h	h�e]r,[  (hh�eeee]r-[  (hheeej [  j [  j [  j [  j [  j [  j [  j [  j [  ]r.[  (jYF  ]r/[  (j[F  ]r0[  (j]F  ]r1[  (h	j�  e]r2[  (hh�e]r3[  (hhe]r4[  (jdF  ]r5[  (h	he]r6[  (hh�e]r7[  (hhe]r8[  (j2R  ]r9[  (h	h�e]r:[  (hh�eeee]r;[  (hheeej.[  ]r<[  (jYF  ]r=[  (j[F  ]r>[  (j]F  ]r?[  (h	j�  e]r@[  (hh�e]rA[  (hhe]rB[  (jdF  ]rC[  (h	he]rD[  (hh�e]rE[  (hhe]rF[  (j2R  ]rG[  (h	h�e]rH[  (hh�eeee]rI[  (hheee]rJ[  (jYF  ]rK[  (j[F  ]rL[  (j]F  ]rM[  (h	j�  e]rN[  (hh�e]rO[  (hhe]rP[  (jdF  ]rQ[  (h	he]rR[  (hh�e]rS[  (hhe]rT[  (j2R  ]rU[  (h	h�e]rV[  (hh�eeee]rW[  (hheeejJ[  ]rX[  (jYF  ]rY[  (j[F  ]rZ[  (j]F  ]r[[  (h	h�e]r\[  (hh�e]r][  (hhe]r^[  (jdF  ]r_[  (h	he]r`[  (hh�e]ra[  (hhe]rb[  (j2R  ]rc[  (h	h�e]rd[  (hh�eeee]re[  (hheeejX[  jX[  jX[  jX[  jX[  ]rf[  (jYF  ]rg[  (j[F  ]rh[  (j]F  ]ri[  (h	h�e]rj[  (hh�e]rk[  (hhe]rl[  (jdF  ]rm[  (h	he]rn[  (hh�e]ro[  (hhe]rp[  (j2R  ]rq[  (h	h�e]rr[  (hh�eeee]rs[  (hheeejf[  jf[  ]rt[  (jYF  ]ru[  (j[F  ]rv[  (j]F  ]rw[  (h	h�e]rx[  (hh�e]ry[  (hhe]rz[  (jdF  ]r{[  (h	he]r|[  (hh�e]r}[  (hhe]r~[  (j2R  ]r[  (h	h�e]r�[  (hh�eeee]r�[  (hheeejt[  jt[  jt[  jt[  ]r�[  (jYF  ]r�[  (j[F  ]r�[  (j]F  ]r�[  (h	h�e]r�[  (hh�e]r�[  (hhe]r�[  (jdF  ]r�[  (h	he]r�[  (hh�e]r�[  (hhe]r�[  (j2R  ]r�[  (h	h�e]r�[  (hh�eeee]r�[  (hheee]r�[  (jYF  ]r�[  (j[F  ]r�[  (j]F  ]r�[  (h	h�e]r�[  (hh�e]r�[  (hhe]r�[  (jdF  ]r�[  (h	he]r�[  (hh�e]r�[  (hhe]r�[  (j2R  ]r�[  (h	h�e]r�[  (hh�eeee]r�[  (hheeej�[  j�[  j�[  ]r�[  (jYF  ]r�[  (j[F  ]r�[  (j]F  ]r�[  (h	h�e]r�[  (hh�e]r�[  (hhe]r�[  (jdF  ]r�[  (h	he]r�[  (hh�e]r�[  (hhe]r�[  (j2R  ]r�[  (h	h�e]r�[  (hh�eeee]r�[  (hheeej�[  ]r�[  (jYF  ]r�[  (j[F  ]r�[  (j]F  ]r�[  (h	h�e]r�[  (hh�e]r�[  (hhe]r�[  (jdF  ]r�[  (h	he]r�[  (hh�e]r�[  (hhe]r�[  (j2R  ]r�[  (h	h�e]r�[  (hh�eeee]r�[  (hheeej�[  ]r�[  (jYF  ]r�[  (j[F  ]r�[  (j]F  ]r�[  (h	j�  e]r�[  (hh�e]r�[  (hhe]r�[  (jdF  ]r�[  (h	he]r�[  (hh�e]r�[  (hhe]r�[  (j2R  ]r�[  (h	h�e]r�[  (hh�eeee]r�[  (hheeej�[  j�[  j�[  j�[  j�[  j�[  j�[  j�[  j�[  j�[  j�[  ]r�[  (jYF  ]r�[  (j[F  ]r�[  (j]F  ]r�[  (h	h�e]r�[  (hh�e]r�[  (hhe]r�[  (jdF  ]r�[  (h	he]r�[  (hh�e]r�[  (hhe]r�[  (j2R  ]r�[  (h	h�e]r�[  (hh�eeee]r�[  (hheeej�[  j�[  j�[  ]r�[  (jYF  ]r�[  (j[F  ]r�[  (j]F  ]r�[  (h	h�e]r�[  (hh�e]r�[  (hhe]r�[  (jdF  ]r�[  (h	he]r�[  (hh�e]r�[  (hhe]r�[  (j2R  ]r�[  (h	h�e]r�[  (hh�eeee]r�[  (hheeej�[  j�[  j�[  j�[  j�[  j�[  j�[  j�[  ]r�[  (jYF  ]r�[  (j[F  ]r�[  (j]F  ]r�[  (h	h�e]r�[  (hh�e]r�[  (hhe]r�[  (jdF  ]r�[  (h	he]r�[  (hh�e]r�[  (hhe]r�[  (j2R  ]r�[  (h	h�e]r�[  (hh�eeee]r�[  (hheeej�[  j�[  j�[  ]r�[  (jYF  ]r�[  (j[F  ]r�[  (j]F  ]r�[  (h	h�e]r�[  (hh�e]r�[  (hhe]r�[  (jdF  ]r�[  (h	he]r�[  (hh�e]r�[  (hhe]r�[  (j2R  ]r�[  (h	h�e]r�[  (hh�eeee]r�[  (hheeej�[  j�[  j�[  j�[  j�[  ]r \  (jYF  ]r\  (j[F  ]r\  (j]F  ]r\  (h	h�e]r\  (hh�e]r\  (hhe]r\  (jdF  ]r\  (h	he]r\  (hh�e]r	\  (hhe]r
\  (j2R  ]r\  (h	h�e]r\  (hh�eeee]r\  (hheeej \  ]r\  (jYF  ]r\  (j[F  ]r\  (j]F  ]r\  (h	h�e]r\  (hh�e]r\  (hhe]r\  (jdF  ]r\  (h	he]r\  (hh�e]r\  (hhe]r\  (j2R  ]r\  (h	h�e]r\  (hh�eeee]r\  (hheeej\  j\  j\  ]r\  (jYF  ]r\  (j[F  ]r\  (j]F  ]r\  (h	h�e]r \  (hh�e]r!\  (hhe]r"\  (jdF  ]r#\  (h	he]r$\  (hh�e]r%\  (hhe]r&\  (j2R  ]r'\  (h	h�e]r(\  (hh�eeee]r)\  (hheeej\  ]r*\  (jYF  ]r+\  (j[F  ]r,\  (j]F  ]r-\  (h	j�  e]r.\  (hh�e]r/\  (hhe]r0\  (jdF  ]r1\  (h	he]r2\  (hh�e]r3\  (hhe]r4\  (j2R  ]r5\  (h	h�e]r6\  (hh�eeee]r7\  (hheeej*\  j*\  j*\  j*\  j*\  j*\  ]r8\  (jYF  ]r9\  (j[F  ]r:\  (j]F  ]r;\  (h	j�  e]r<\  (hh�e]r=\  (hhe]r>\  (jdF  ]r?\  (h	he]r@\  (hh�e]rA\  (hhe]rB\  (j2R  ]rC\  (h	h�e]rD\  (hh�eeee]rE\  (hheeej8\  j8\  j8\  j8\  j8\  j8\  j8\  j8\  ]rF\  (jYF  ]rG\  (j[F  ]rH\  (j]F  ]rI\  (h	j�  e]rJ\  (hh�e]rK\  (hhe]rL\  (jdF  ]rM\  (h	he]rN\  (hh�e]rO\  (hhe]rP\  (j2R  ]rQ\  (h	h�e]rR\  (hh�eeee]rS\  (hheeejF\  jF\  jF\  jF\  jF\  jF\  jF\  jF\  jF\  jF\  jF\  jF\  jF\  jF\  ]rT\  (jYF  ]rU\  (j[F  ]rV\  (j]F  ]rW\  (h	j�  e]rX\  (hh�e]rY\  (hhe]rZ\  (jdF  ]r[\  (h	he]r\\  (hh�e]r]\  (hhe]r^\  (j2R  ]r_\  (h	h�e]r`\  (hh�eeee]ra\  (hheeejT\  jT\  ]rb\  (jYF  ]rc\  (j[F  ]rd\  (j]F  ]re\  (h	j�  e]rf\  (hh�e]rg\  (hhe]rh\  (jdF  ]ri\  (h	he]rj\  (hh�e]rk\  (hhe]rl\  (j2R  ]rm\  (h	h�e]rn\  (hh�eeee]ro\  (hheeejb\  jb\  jb\  ]rp\  (jYF  ]rq\  (j[F  ]rr\  (j]F  ]rs\  (h	j�  e]rt\  (hh�e]ru\  (hhe]rv\  (jdF  ]rw\  (h	he]rx\  (hh�e]ry\  (hhe]rz\  (j2R  ]r{\  (h	h�e]r|\  (hh�eeee]r}\  (hheeejp\  jp\  jp\  jp\  jp\  ]r~\  (jYF  ]r\  (j[F  ]r�\  (j]F  ]r�\  (h	j�  e]r�\  (hh�e]r�\  (hhe]r�\  (jdF  ]r�\  (h	he]r�\  (hh�e]r�\  (hhe]r�\  (j2R  ]r�\  (h	h�e]r�\  (hh�eeee]r�\  (hheeej~\  j~\  j~\  j~\  j~\  j~\  j~\  j~\  j~\  ]r�\  (jYF  ]r�\  (j[F  ]r�\  (j]F  ]r�\  (h	j�  e]r�\  (hh�e]r�\  (hhe]r�\  (jdF  ]r�\  (h	he]r�\  (hh�e]r�\  (hhe]r�\  (j2R  ]r�\  (h	h�e]r�\  (hh�eeee]r�\  (hheeej�\  j�\  ]r�\  (jYF  ]r�\  (j[F  ]r�\  (j]F  ]r�\  (h	j�  e]r�\  (hh�e]r�\  (hhe]r�\  (jdF  ]r�\  (h	he]r�\  (hh�e]r�\  (hhe]r�\  (j2R  ]r�\  (h	h�e]r�\  (hh�eeee]r�\  (hheeej�\  ]r�\  (jYF  ]r�\  (j[F  ]r�\  (j]F  ]r�\  (h	j�  e]r�\  (hh�e]r�\  (hhe]r�\  (jdF  ]r�\  (h	he]r�\  (hh�e]r�\  (hhe]r�\  (j2R  ]r�\  (h	h�e]r�\  (hh�eeee]r�\  (hheeej�\  j�\  j�\  ]r�\  (jYF  ]r�\  (j[F  ]r�\  (j]F  ]r�\  (h	j�  e]r�\  (hh�e]r�\  (hhe]r�\  (jdF  ]r�\  (h	he]r�\  (hh�e]r�\  (hhe]r�\  (j2R  ]r�\  (h	h�e]r�\  (hh�eeee]r�\  (hheeej�\  j�\  ]r�\  (jYF  ]r�\  (j[F  ]r�\  (j]F  ]r�\  (h	j�  e]r�\  (hh�e]r�\  (hhe]r�\  (jdF  ]r�\  (h	he]r�\  (hh�e]r�\  (hhe]r�\  (j2R  ]r�\  (h	h�e]r�\  (hh�eeee]r�\  (hheeej�\  j�\  ]r�\  (jYF  ]r�\  (j[F  ]r�\  (j]F  ]r�\  (h	j�  e]r�\  (hh�e]r�\  (hhe]r�\  (jdF  ]r�\  (h	he]r�\  (hh�e]r�\  (hhe]r�\  (j2R  ]r�\  (h	h�e]r�\  (hh�eeee]r�\  (hheeej�\  j�\  j�\  j�\  j�\  j�\  j�\  ]r�\  (jYF  ]r�\  (j[F  ]r�\  (j]F  ]r�\  (h	j�  e]r�\  (hh�e]r�\  (hhe]r�\  (jdF  ]r�\  (h	he]r�\  (hh�e]r�\  (hhe]r�\  (j2R  ]r�\  (h	h�e]r�\  (hh�eeee]r�\  (hheeej�\  j�\  j�\  j�\  ]r�\  (jYF  ]r�\  (j[F  ]r�\  (j]F  ]r�\  (h	j�  e]r�\  (hh�e]r�\  (hhe]r�\  (jdF  ]r�\  (h	he]r�\  (hh�e]r�\  (hhe]r�\  (j2R  ]r�\  (h	h�e]r�\  (hh�eeee]r�\  (hheeej�\  ]r�\  (jYF  ]r�\  (j[F  ]r�\  (j]F  ]r�\  (h	j�  e]r ]  (hh�e]r]  (hhe]r]  (jdF  ]r]  (h	he]r]  (hh�e]r]  (hhe]r]  (j2R  ]r]  (h	h�e]r]  (hh�eeee]r	]  (hheeej�\  j�\  j�\  j�\  j�\  j�\  j�\  j�\  j�\  j�\  j�\  j�\  j�\  ]r
]  (jYF  ]r]  (j[F  ]r]  (j]F  ]r]  (h	j�  e]r]  (hh�e]r]  (hhe]r]  (jdF  ]r]  (h	he]r]  (hh�e]r]  (hhe]r]  (j2R  ]r]  (h	h�e]r]  (hh�eeee]r]  (hheeej
]  j
]  j
]  j
]  j
]  j
]  j
]  j
]  j
]  j
]  j
]  j
]  ]r]  (jYF  ]r]  (j[F  ]r]  (j]F  ]r]  (h	j�  e]r]  (hh�e]r]  (hhe]r]  (jdF  ]r]  (h	he]r ]  (hh�e]r!]  (hhe]r"]  (j2R  ]r#]  (h	h�e]r$]  (hh�eeee]r%]  (hheeej]  j]  j]  j]  j]  j]  j]  j]  j]  j]  j]  j]  j]  j]  ]r&]  (jYF  ]r']  (j[F  ]r(]  (j]F  ]r)]  (h	j�  e]r*]  (hh�e]r+]  (hhe]r,]  (jdF  ]r-]  (h	he]r.]  (hh�e]r/]  (hhe]r0]  (j2R  ]r1]  (h	h�e]r2]  (hh�eeee]r3]  (hheeej&]  j&]  ]r4]  (jYF  ]r5]  (j[F  ]r6]  (j]F  ]r7]  (h	j�  e]r8]  (hh�e]r9]  (hhe]r:]  (jdF  ]r;]  (h	he]r<]  (hh�e]r=]  (hhe]r>]  (j2R  ]r?]  (h	h�e]r@]  (hh�eeee]rA]  (hheeej4]  ]rB]  (jYF  ]rC]  (j[F  ]rD]  (j]F  ]rE]  (h	j�  e]rF]  (hh�e]rG]  (hhe]rH]  (jdF  ]rI]  (h	he]rJ]  (hh�e]rK]  (hhe]rL]  (j2R  ]rM]  (h	h�e]rN]  (hh�eeee]rO]  (hheeejB]  jB]  jB]  jB]  jB]  jB]  ]rP]  (jYF  ]rQ]  (j[F  ]rR]  (j]F  ]rS]  (h	j�  e]rT]  (hh�e]rU]  (hhe]rV]  (jdF  ]rW]  (h	he]rX]  (hh�e]rY]  (hhe]rZ]  (j2R  ]r[]  (h	h�e]r\]  (hh�eeee]r]]  (hheeejP]  ]r^]  (jYF  ]r_]  (j[F  ]r`]  (j]F  ]ra]  (h	j�  e]rb]  (hh�e]rc]  (hhe]rd]  (jdF  ]re]  (h	he]rf]  (hh�e]rg]  (hhe]rh]  (j2R  ]ri]  (h	h�e]rj]  (hh�eeee]rk]  (hheeej^]  j^]  j^]  j^]  j^]  j^]  j^]  j^]  ]rl]  (jYF  ]rm]  (j[F  ]rn]  (j]F  ]ro]  (h	j�  e]rp]  (hh�e]rq]  (hhe]rr]  (jdF  ]rs]  (h	he]rt]  (hh�e]ru]  (hhe]rv]  (j2R  ]rw]  (h	h�e]rx]  (hh�eeee]ry]  (hheee]rz]  (jYF  ]r{]  (j[F  ]r|]  (j]F  ]r}]  (h	j�  e]r~]  (hh�e]r]  (hhe]r�]  (jdF  ]r�]  (h	he]r�]  (hh�e]r�]  (hhe]r�]  (j2R  ]r�]  (h	h�e]r�]  (hh�eeee]r�]  (hheeejz]  jz]  jz]  jz]  jz]  jz]  ]r�]  (jYF  ]r�]  (j[F  ]r�]  (j]F  ]r�]  (h	j�  e]r�]  (hh�e]r�]  (hhe]r�]  (jdF  ]r�]  (h	he]r�]  (hh�e]r�]  (hhe]r�]  (j2R  ]r�]  (h	h�e]r�]  (hh�eeee]r�]  (hheeej�]  j�]  j�]  j�]  j�]  j�]  j�]  j�]  j�]  ]r�]  (jYF  ]r�]  (j[F  ]r�]  (j]F  ]r�]  (h	j�  e]r�]  (hh�e]r�]  (hhe]r�]  (jdF  ]r�]  (h	he]r�]  (hh�e]r�]  (hhe]r�]  (j2R  ]r�]  (h	h�e]r�]  (hh�eeee]r�]  (hheeej�]  j�]  j�]  ]r�]  (jYF  ]r�]  (j[F  ]r�]  (j]F  ]r�]  (h	j�  e]r�]  (hh�e]r�]  (hhe]r�]  (jdF  ]r�]  (h	he]r�]  (hh�e]r�]  (hhe]r�]  (j2R  ]r�]  (h	h�e]r�]  (hh�eeee]r�]  (hheeej�]  j�]  j�]  j�]  ]r�]  (jYF  ]r�]  (j[F  ]r�]  (j]F  ]r�]  (h	j�  e]r�]  (hh�e]r�]  (hhe]r�]  (jdF  ]r�]  (h	he]r�]  (hh�e]r�]  (hhe]r�]  (j2R  ]r�]  (h	h�e]r�]  (hh�eeee]r�]  (hheeej�]  j�]  j�]  ]r�]  (jYF  ]r�]  (j[F  ]r�]  (j]F  ]r�]  (h	j�  e]r�]  (hh�e]r�]  (hhe]r�]  (jdF  ]r�]  (h	he]r�]  (hh�e]r�]  (hhe]r�]  (j2R  ]r�]  (h	h�e]r�]  (hh�eeee]r�]  (hheeej�]  j�]  j�]  j�]  j�]  j�]  j�]  j�]  j�]  j�]  ]r�]  (jYF  ]r�]  (j[F  ]r�]  (j]F  ]r�]  (h	j�  e]r�]  (hh�e]r�]  (hhe]r�]  (jdF  ]r�]  (h	he]r�]  (hh�e]r�]  (hhe]r�]  (j2R  ]r�]  (h	h�e]r�]  (hh�eeee]r�]  (hheeej�]  j�]  j�]  ]r�]  (jYF  ]r�]  (j[F  ]r�]  (j]F  ]r�]  (h	j�  e]r�]  (hh�e]r�]  (hhe]r�]  (jdF  ]r�]  (h	he]r�]  (hh�e]r�]  (hhe]r�]  (j2R  ]r�]  (h	h�e]r�]  (hh�eeee]r�]  (hheee]r�]  (jYF  ]r�]  (j[F  ]r�]  (j]F  ]r�]  (h	j�  e]r�]  (hh�e]r�]  (hhe]r�]  (jdF  ]r�]  (h	he]r�]  (hh�e]r�]  (hhe]r�]  (j2R  ]r�]  (h	h�e]r�]  (hh�eeee]r�]  (hheeej�]  j�]  ]r�]  (jYF  ]r�]  (j[F  ]r�]  (j]F  ]r�]  (h	j�  e]r�]  (hh�e]r�]  (hhe]r�]  (jdF  ]r�]  (h	he]r ^  (hh�e]r^  (hhe]r^  (j2R  ]r^  (h	h�e]r^  (hh�eeee]r^  (hheeej�]  j�]  j�]  ]r^  (jYF  ]r^  (j[F  ]r^  (j]F  ]r	^  (h	j�  e]r
^  (hh�e]r^  (hhe]r^  (jdF  ]r^  (h	he]r^  (hh�e]r^  (hhe]r^  (j2R  ]r^  (h	h�e]r^  (hh�eeee]r^  (hheeej^  j^  j^  j^  j^  j^  j^  ]r^  (jYF  ]r^  (X   Oblr^  ]r^  (jD>  ]r^  (h	h�e]r^  (hh�e]r^  (hhe]r^  (jD>  ]r^  (h	h
e]r^  (hh<e]r^  (hhe]r^  (X	   Next-Mover ^  ]r!^  (h	he]r"^  (hh�eeee]r#^  (hheee]r$^  (jYF  ]r%^  (j^  ]r&^  (jD>  ]r'^  (h	h�e]r(^  (hh�e]r)^  (hhe]r*^  (jD>  ]r+^  (h	h
e]r,^  (hh<e]r-^  (hhe]r.^  (j ^  ]r/^  (h	he]r0^  (hh�eeee]r1^  (hheeej$^  j$^  j$^  j$^  ]r2^  (jYF  ]r3^  (j^  ]r4^  (jD>  ]r5^  (h	h�e]r6^  (hh�e]r7^  (hhe]r8^  (jD>  ]r9^  (h	h
e]r:^  (hh�e]r;^  (hhe]r<^  (j ^  ]r=^  (h	he]r>^  (hh�eeee]r?^  (hheeej2^  ]r@^  (jYF  ]rA^  (j^  ]rB^  (jD>  ]rC^  (h	h�e]rD^  (hh�e]rE^  (hhe]rF^  (jD>  ]rG^  (h	h�e]rH^  (hh�e]rI^  (hhe]rJ^  (j ^  ]rK^  (h	he]rL^  (hh�eeee]rM^  (hheeej@^  j@^  j@^  ]rN^  (jYF  ]rO^  (j^  ]rP^  (jD>  ]rQ^  (h	h�e]rR^  (hh�e]rS^  (hhe]rT^  (jD>  ]rU^  (h	h�e]rV^  (hh�e]rW^  (hhe]rX^  (j ^  ]rY^  (h	he]rZ^  (hh�eeee]r[^  (hheeejN^  jN^  jN^  jN^  jN^  jN^  jN^  ]r\^  (jYF  ]r]^  (j^  ]r^^  (jD>  ]r_^  (h	h�e]r`^  (hh�e]ra^  (hhe]rb^  (jD>  ]rc^  (h	h�e]rd^  (hh�e]re^  (hhe]rf^  (j ^  ]rg^  (h	he]rh^  (hh�eeee]ri^  (hheee]rj^  (jYF  ]rk^  (j^  ]rl^  (jD>  ]rm^  (h	h�e]rn^  (hh�e]ro^  (hhe]rp^  (jD>  ]rq^  (h	h�e]rr^  (hh�e]rs^  (hhe]rt^  (j ^  ]ru^  (h	he]rv^  (hh�eeee]rw^  (hheeejj^  jj^  jj^  jj^  jj^  jj^  ]rx^  (jYF  ]ry^  (j^  ]rz^  (jD>  ]r{^  (h	h�e]r|^  (hh�e]r}^  (hhe]r~^  (jD>  ]r^  (h	h�e]r�^  (hh�e]r�^  (hhe]r�^  (j ^  ]r�^  (h	he]r�^  (hh�eeee]r�^  (hheeejx^  jx^  jx^  jx^  jx^  jx^  jx^  ]r�^  (jYF  ]r�^  (j^  ]r�^  (jD>  ]r�^  (h	h�e]r�^  (hh�e]r�^  (hhe]r�^  (jD>  ]r�^  (h	h�e]r�^  (hh�e]r�^  (hhe]r�^  (j ^  ]r�^  (h	he]r�^  (hh�eeee]r�^  (hheeej�^  ]r�^  (jYF  ]r�^  (j^  ]r�^  (jD>  ]r�^  (h	h�e]r�^  (hh�e]r�^  (hhe]r�^  (jD>  ]r�^  (h	h�e]r�^  (hh�e]r�^  (hhe]r�^  (j ^  ]r�^  (h	he]r�^  (hh�eeee]r�^  (hheeej�^  j�^  j�^  j�^  ]r�^  (jYF  ]r�^  (j^  ]r�^  (jD>  ]r�^  (h	h�e]r�^  (hh�e]r�^  (hhe]r�^  (jD>  ]r�^  (h	h�e]r�^  (hh�e]r�^  (hhe]r�^  (j ^  ]r�^  (h	he]r�^  (hh�eeee]r�^  (hheeej�^  j�^  ]r�^  (jYF  ]r�^  (j^  ]r�^  (jD>  ]r�^  (h	h�e]r�^  (hh�e]r�^  (hhe]r�^  (jD>  ]r�^  (h	h�e]r�^  (hh�e]r�^  (hhe]r�^  (j ^  ]r�^  (h	he]r�^  (hh�eeee]r�^  (hheeej�^  j�^  j�^  j�^  e(j�^  e]r�^  (]r�^  (X   Normsr�^  ]r�^  (X   Oblr�^  ]r�^  (X   Movedr�^  ]r�^  (h	he]r�^  (hX   anyr�^  e]r�^  (hhe]r�^  (X   Movedr�^  ]r�^  (h	X   anyr�^  e]r�^  (hX   triangler�^  e]r�^  (hhe]r�^  (X	   Next-Mover�^  ]r�^  (h	X   anyr�^  e]r�^  (hX   anyr�^  eeee]r�^  (hhee]r�^  (h!]r�^  (h#h$e]r�^  (h	X   anyr�^  e]r�^  (hX   squarer�^  e]r�^  (h)X   anyr�^  eeej�^  ]r�^  (j�^  ]r�^  (j�^  ]r�^  (j�^  ]r�^  (h	he]r�^  (hj�^  e]r�^  (hhe]r�^  (j�^  ]r�^  (h	j�^  e]r�^  (hj�^  e]r�^  (hhe]r�^  (j�^  ]r�^  (h	j�^  e]r�^  (hj�^  eeee]r�^  (hhee]r�^  (h!]r�^  (h#h$e]r�^  (h	j�^  e]r�^  (hj�^  e]r�^  (h)heeej�^  j�^  ]r�^  (j�^  ]r�^  (j�^  ]r�^  (j�^  ]r�^  (h	he]r�^  (hj�^  e]r�^  (hhe]r�^  (j�^  ]r�^  (h	j�^  e]r�^  (hj�^  e]r�^  (hhe]r�^  (j�^  ]r�^  (h	j�^  e]r�^  (hj�^  eeee]r�^  (hhee]r _  (h!]r_  (h#h$e]r_  (h	j�  e]r_  (hh�e]r_  (h)h�eee]r_  (j�^  ]r_  (j�^  ]r_  (j�^  ]r_  (h	he]r	_  (hj�^  e]r
_  (hhe]r_  (j�^  ]r_  (h	j�^  e]r_  (hj�^  e]r_  (hhe]r_  (j�^  ]r_  (h	j�^  e]r_  (hj�^  eeee]r_  (hhee]r_  (h!]r_  (h#h$e]r_  (h	j�  e]r_  (hh�e]r_  (h)h�eeej_  ]r_  (j�^  ]r_  (j�^  ]r_  (j�^  ]r_  (h	he]r_  (hj�^  e]r_  (hhe]r_  (j�^  ]r_  (h	j�^  e]r _  (hj�^  e]r!_  (hhe]r"_  (j�^  ]r#_  (h	j�^  e]r$_  (hj�^  eeee]r%_  (hhee]r&_  (h!]r'_  (h#h$e]r(_  (h	j�  e]r)_  (hh�e]r*_  (h)h�eeej_  j_  ]r+_  (j�^  ]r,_  (j�^  ]r-_  (j�^  ]r._  (h	he]r/_  (hj�^  e]r0_  (hhe]r1_  (j�^  ]r2_  (h	j�^  e]r3_  (hj�^  e]r4_  (hhe]r5_  (j�^  ]r6_  (h	j�^  e]r7_  (hj�^  eeee]r8_  (hhee]r9_  (h!]r:_  (h#h$e]r;_  (h	j�  e]r<_  (hh�e]r=_  (h)heeej+_  j+_  ]r>_  (j�^  ]r?_  (j�^  ]r@_  (j�^  ]rA_  (h	he]rB_  (hj�^  e]rC_  (hhe]rD_  (j�^  ]rE_  (h	j�^  e]rF_  (hj�^  e]rG_  (hhe]rH_  (j�^  ]rI_  (h	j�^  e]rJ_  (hj�^  eeee]rK_  (hhee]rL_  (h!]rM_  (h#h$e]rN_  (h	j�  e]rO_  (hh�e]rP_  (h)heee]rQ_  (j�^  ]rR_  (j�^  ]rS_  (j�^  ]rT_  (h	he]rU_  (hj�^  e]rV_  (hhe]rW_  (j�^  ]rX_  (h	j�^  e]rY_  (hj�^  e]rZ_  (hhe]r[_  (j�^  ]r\_  (h	j�^  e]r]_  (hj�^  eeee]r^_  (hhee]r__  (h!]r`_  (h#h$e]ra_  (h	j�  e]rb_  (hh�e]rc_  (h)heee]rd_  (j�^  ]re_  (j�^  ]rf_  (j�^  ]rg_  (h	he]rh_  (hj�^  e]ri_  (hhe]rj_  (j�^  ]rk_  (h	j�^  e]rl_  (hj�^  e]rm_  (hhe]rn_  (j�^  ]ro_  (h	j�^  e]rp_  (hj�^  eeee]rq_  (hhee]rr_  (h!]rs_  (h#h$e]rt_  (h	j�  e]ru_  (hh�e]rv_  (h)heeejd_  ]rw_  (j�^  ]rx_  (j�^  ]ry_  (j�^  ]rz_  (h	he]r{_  (hj�^  e]r|_  (hhe]r}_  (j�^  ]r~_  (h	j�^  e]r_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hj�^  eeee]r�_  (hhee]r�_  (h!]r�_  (h#h$e]r�_  (h	j�  e]r�_  (hh�e]r�_  (h)heeejw_  jw_  ]r�_  (j�^  ]r�_  (j�^  ]r�_  (j�^  ]r�_  (h	he]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hj�^  eeee]r�_  (hhee]r�_  (h!]r�_  (h#h$e]r�_  (h	j�  e]r�_  (hh�e]r�_  (h)heee]r�_  (j�^  ]r�_  (j�^  ]r�_  (j�^  ]r�_  (h	he]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hh<eeee]r�_  (hhee]r�_  (h!]r�_  (h#h$e]r�_  (h	j�  e]r�_  (hh�e]r�_  (h)heee]r�_  (j�^  ]r�_  (j�^  ]r�_  (j�^  ]r�_  (h	he]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hh<eeee]r�_  (hhee]r�_  (h!]r�_  (h#h$e]r�_  (h	j�  e]r�_  (hh�e]r�_  (h)heeej�_  ]r�_  (j�^  ]r�_  (j�^  ]r�_  (j�^  ]r�_  (h	he]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hh<eeee]r�_  (hhee]r�_  (h!]r�_  (h#h$e]r�_  (h	j�  e]r�_  (hh<e]r�_  (h)heeej�_  ]r�_  (j�^  ]r�_  (j�^  ]r�_  (j�^  ]r�_  (h	he]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hh<eeee]r�_  (hhee]r�_  (h!]r�_  (h#h$e]r�_  (h	j�  e]r�_  (hh<e]r�_  (h)heeej�_  j�_  ]r�_  (j�^  ]r�_  (j�^  ]r�_  (j�^  ]r�_  (h	he]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hj�^  e]r�_  (hhe]r�_  (j�^  ]r�_  (h	j�^  e]r�_  (hh<eeee]r�_  (hhee]r�_  (h!]r�_  (h#h$e]r�_  (h	j�  e]r�_  (hh<e]r�_  (h)heee]r�_  (j�^  ]r�_  (j�^  ]r�_  (j�^  ]r�_  (h	h�e]r `  (hj�^  e]r`  (hhe]r`  (j�^  ]r`  (h	j�^  e]r`  (hj�^  e]r`  (hhe]r`  (j�^  ]r`  (h	j�^  e]r`  (hh<eeee]r	`  (hhee]r
`  (h!]r`  (h#h$e]r`  (h	j�  e]r`  (hh<e]r`  (h)heee]r`  (j�^  ]r`  (j�^  ]r`  (j�^  ]r`  (h	h�e]r`  (hj�^  e]r`  (hhe]r`  (j�^  ]r`  (h	j�^  e]r`  (hj�^  e]r`  (hhe]r`  (j�^  ]r`  (h	j�^  e]r`  (hh<eeee]r`  (hhee]r`  (h!]r`  (h#h$e]r`  (h	j�  e]r `  (hh<e]r!`  (h)heee]r"`  (j�^  ]r#`  (j�^  ]r$`  (j�^  ]r%`  (h	h�e]r&`  (hj�^  e]r'`  (hhe]r(`  (j�^  ]r)`  (h	j�^  e]r*`  (hj�^  e]r+`  (hhe]r,`  (j�^  ]r-`  (h	j�^  e]r.`  (hh<eeee]r/`  (hhee]r0`  (h!]r1`  (h#h$e]r2`  (h	j�  e]r3`  (hh<e]r4`  (h)heeej"`  ]r5`  (j�^  ]r6`  (j�^  ]r7`  (j�^  ]r8`  (h	h�e]r9`  (hj�^  e]r:`  (hhe]r;`  (j�^  ]r<`  (h	he]r=`  (hj�^  e]r>`  (hhe]r?`  (j�^  ]r@`  (h	j�^  e]rA`  (hh<eeee]rB`  (hhee]rC`  (h!]rD`  (h#h$e]rE`  (h	j�  e]rF`  (hh<e]rG`  (h)heeej5`  j5`  j5`  j5`  j5`  j5`  ]rH`  (j�^  ]rI`  (j�^  ]rJ`  (j�^  ]rK`  (h	h�e]rL`  (hj�^  e]rM`  (hhe]rN`  (j�^  ]rO`  (h	he]rP`  (hj�^  e]rQ`  (hhe]rR`  (j�^  ]rS`  (h	j�^  e]rT`  (hh<eeee]rU`  (hhee]rV`  (h!]rW`  (h#h$e]rX`  (h	he]rY`  (hh<e]rZ`  (h)heeejH`  jH`  ]r[`  (j�^  ]r\`  (j�^  ]r]`  (j�^  ]r^`  (h	h�e]r_`  (hj�^  e]r``  (hhe]ra`  (j�^  ]rb`  (h	he]rc`  (hj�^  e]rd`  (hhe]re`  (j�^  ]rf`  (h	j�^  e]rg`  (hh<eeee]rh`  (hhee]ri`  (h!]rj`  (h#h$e]rk`  (h	he]rl`  (hh<e]rm`  (h)heeej[`  j[`  j[`  ]rn`  (j�^  ]ro`  (j�^  ]rp`  (j�^  ]rq`  (h	h�e]rr`  (hj�^  e]rs`  (hhe]rt`  (j�^  ]ru`  (h	he]rv`  (hj�^  e]rw`  (hhe]rx`  (j�^  ]ry`  (h	j�^  e]rz`  (hh<eeee]r{`  (hhee]r|`  (h!]r}`  (h#h$e]r~`  (h	he]r`  (hh�e]r�`  (h)heeejn`  jn`  jn`  jn`  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (h	h�e]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	he]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	j�^  e]r�`  (hh<eeee]r�`  (hhee]r�`  (h!]r�`  (h#h$e]r�`  (h	he]r�`  (hh�e]r�`  (h)heee]r�`  (j�^  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (h	h�e]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	he]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	j�^  e]r�`  (hh<eeee]r�`  (hhee]r�`  (h!]r�`  (h#h$e]r�`  (h	h
e]r�`  (hh�e]r�`  (h)heeej�`  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (h	h�e]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	he]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	j�^  e]r�`  (hh<eeee]r�`  (hhee]r�`  (h!]r�`  (h#h$e]r�`  (h	h
e]r�`  (hh�e]r�`  (h)heeej�`  j�`  j�`  j�`  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (h	h�e]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	h�e]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	j�^  e]r�`  (hh<eeee]r�`  (hhee]r�`  (h!]r�`  (h#h$e]r�`  (h	h
e]r�`  (hh�e]r�`  (h)heee]r�`  (j�^  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (h	h�e]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	h�e]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	j�^  e]r�`  (hh<eeee]r�`  (hhee]r�`  (h!]r�`  (h#h$e]r�`  (h	he]r�`  (hh�e]r�`  (h)heeej�`  j�`  j�`  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (h	h�e]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	h�e]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	j�^  e]r�`  (hh<eeee]r�`  (hhee]r�`  (h!]r�`  (h#h$e]r�`  (h	j�  e]r�`  (hh�e]r�`  (h)heeej�`  j�`  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (j�^  ]r�`  (h	h�e]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	h�e]r�`  (hj�^  e]r�`  (hhe]r�`  (j�^  ]r�`  (h	j�^  e]r�`  (hh<eeee]r a  (hhee]ra  (h!]ra  (h#h$e]ra  (h	j�  e]ra  (hh�e]ra  (h)heeej�`  j�`  ]ra  (j�^  ]ra  (j�^  ]ra  (j�^  ]r	a  (h	h�e]r
a  (hj�^  e]ra  (hhe]ra  (j�^  ]ra  (h	h�e]ra  (hj�^  e]ra  (hhe]ra  (j�^  ]ra  (h	j�^  e]ra  (hh<eeee]ra  (hhee]ra  (h!]ra  (h#h$e]ra  (h	j�  e]ra  (hh�e]ra  (h)heee]ra  (j�^  ]ra  (j�^  ]ra  (j�^  ]ra  (h	h�e]ra  (hj�^  e]ra  (hhe]ra  (j�^  ]r a  (h	h�e]r!a  (hj�^  e]r"a  (hhe]r#a  (j�^  ]r$a  (h	j�^  e]r%a  (hh<eeee]r&a  (hhee]r'a  (h!]r(a  (h#h$e]r)a  (h	j�  e]r*a  (hh�e]r+a  (h)heee]r,a  (j�^  ]r-a  (j�^  ]r.a  (j�^  ]r/a  (h	h�e]r0a  (hj�^  e]r1a  (hhe]r2a  (j�^  ]r3a  (h	h�e]r4a  (hj�^  e]r5a  (hhe]r6a  (j�^  ]r7a  (h	j�^  e]r8a  (hh<eeee]r9a  (hhee]r:a  (h!]r;a  (h#h$e]r<a  (h	j�  e]r=a  (hh�e]r>a  (h)heee]r?a  (j�^  ]r@a  (j�^  ]rAa  (j�^  ]rBa  (h	h�e]rCa  (hj�^  e]rDa  (hhe]rEa  (j�^  ]rFa  (h	h�e]rGa  (hj�^  e]rHa  (hhe]rIa  (j�^  ]rJa  (h	j�^  e]rKa  (hh<eeee]rLa  (hhee]rMa  (h!]rNa  (h#h$e]rOa  (h	j�  e]rPa  (hh<e]rQa  (h)heee]rRa  (j�^  ]rSa  (j�^  ]rTa  (j�^  ]rUa  (h	h�e]rVa  (hj�^  e]rWa  (hhe]rXa  (j�^  ]rYa  (h	h�e]rZa  (hh�e]r[a  (hhe]r\a  (j�^  ]r]a  (h	j�^  e]r^a  (hh<eeee]r_a  (hhee]r`a  (h!]raa  (h#h$e]rba  (h	j�  e]rca  (hh<e]rda  (h)heeejRa  ]rea  (j�^  ]rfa  (j�^  ]rga  (j�^  ]rha  (h	h�e]ria  (hh�e]rja  (hhe]rka  (j�^  ]rla  (h	h�e]rma  (hh�e]rna  (hhe]roa  (j�^  ]rpa  (h	j�^  e]rqa  (hh<eeee]rra  (hhee]rsa  (h!]rta  (h#h$e]rua  (h	j�  e]rva  (hh<e]rwa  (h)heeejea  jea  jea  jea  ]rxa  (j�^  ]rya  (j�^  ]rza  (j�^  ]r{a  (h	h�e]r|a  (hh�e]r}a  (hhe]r~a  (j�^  ]ra  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	j�^  e]r�a  (hh<eeee]r�a  (hhee]r�a  (h!]r�a  (h#h$e]r�a  (h	j�  e]r�a  (hh<e]r�a  (h)heee]r�a  (j�^  ]r�a  (j�^  ]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	j�^  e]r�a  (hh<eeee]r�a  (hhee]r�a  (h!]r�a  (h#h$e]r�a  (h	j�  e]r�a  (hh<e]r�a  (h)heeej�a  j�a  j�a  j�a  j�a  ]r�a  (j�^  ]r�a  (j�^  ]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	j�^  e]r�a  (hh<eeee]r�a  (hhee]r�a  (h!]r�a  (h#h$e]r�a  (h	j�  e]r�a  (hh<e]r�a  (h)heeej�a  j�a  j�a  ]r�a  (j�^  ]r�a  (j�^  ]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	j�^  e]r�a  (hh<eeee]r�a  (hhee]r�a  (h!]r�a  (h#h$e]r�a  (h	j�  e]r�a  (hh<e]r�a  (h)heeej�a  ]r�a  (j�^  ]r�a  (j�^  ]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	j�^  e]r�a  (hh<eeee]r�a  (hhee]r�a  (h!]r�a  (h#h$e]r�a  (h	j�  e]r�a  (hh<e]r�a  (h)heeej�a  j�a  ]r�a  (j�^  ]r�a  (j�^  ]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	h
e]r�a  (hh<eeee]r�a  (hhee]r�a  (h!]r�a  (h#h$e]r�a  (h	j�  e]r�a  (hh<e]r�a  (h)heeej�a  ]r�a  (j�^  ]r�a  (j�^  ]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	h�e]r�a  (hh�e]r�a  (hhe]r�a  (j�^  ]r�a  (h	h
e]r�a  (hh<eeee]r�a  (hhee]r�a  (h!]r�a  (h#h$e]r�a  (h	j�  e]r�a  (hh<e]r�a  (h)heee]r�a  (j�^  ]r�a  (j�^  ]r�a  (j�^  ]r b  (h	h�e]rb  (hh�e]rb  (hhe]rb  (j�^  ]rb  (h	h�e]rb  (hh�e]rb  (hhe]rb  (j�^  ]rb  (h	h
e]r	b  (hh<eeee]r
b  (hhee]rb  (h!]rb  (h#h$e]rb  (h	j�  e]rb  (hh<e]rb  (h)heee]rb  (j�^  ]rb  (j�^  ]rb  (j�^  ]rb  (h	h�e]rb  (hh�e]rb  (hhe]rb  (j�^  ]rb  (h	h�e]rb  (hh�e]rb  (hhe]rb  (j�^  ]rb  (h	h
e]rb  (hh<eeee]rb  (hhee]rb  (h!]rb  (h#h$e]r b  (h	j�  e]r!b  (hh<e]r"b  (h)heeejb  ]r#b  (j�^  ]r$b  (j�^  ]r%b  (j�^  ]r&b  (h	h�e]r'b  (hh�e]r(b  (hhe]r)b  (j�^  ]r*b  (h	h�e]r+b  (hh�e]r,b  (hhe]r-b  (j�^  ]r.b  (h	h
e]r/b  (hh<eeee]r0b  (hhee]r1b  (h!]r2b  (h#h$e]r3b  (h	j�  e]r4b  (hh<e]r5b  (h)heeej#b  j#b  ]r6b  (j�^  ]r7b  (j�^  ]r8b  (j�^  ]r9b  (h	h�e]r:b  (hh�e]r;b  (hhe]r<b  (j�^  ]r=b  (h	h�e]r>b  (hh�e]r?b  (hhe]r@b  (j�^  ]rAb  (h	h
e]rBb  (hh<eeee]rCb  (hhee]rDb  (h!]rEb  (h#h$e]rFb  (h	j�  e]rGb  (hh<e]rHb  (h)h�eee]rIb  (j�^  ]rJb  (j�^  ]rKb  (j�^  ]rLb  (h	h�e]rMb  (hh�e]rNb  (hhe]rOb  (j�^  ]rPb  (h	h�e]rQb  (hh�e]rRb  (hhe]rSb  (j�^  ]rTb  (h	h
e]rUb  (hh<eeee]rVb  (hhee]rWb  (h!]rXb  (h#h$e]rYb  (h	j�  e]rZb  (hh<e]r[b  (h)h�eee]r\b  (j�^  ]r]b  (j�^  ]r^b  (j�^  ]r_b  (h	h�e]r`b  (hh�e]rab  (hhe]rbb  (j�^  ]rcb  (h	h�e]rdb  (hh�e]reb  (hhe]rfb  (j�^  ]rgb  (h	h
e]rhb  (hh<eeee]rib  (hhee]rjb  (h!]rkb  (h#h$e]rlb  (h	j�  e]rmb  (hh<e]rnb  (h)h�eee]rob  (j�^  ]rpb  (j�^  ]rqb  (j�^  ]rrb  (h	h�e]rsb  (hh�e]rtb  (hhe]rub  (j�^  ]rvb  (h	h�e]rwb  (hh�e]rxb  (hhe]ryb  (j�^  ]rzb  (h	h
e]r{b  (hh<eeee]r|b  (hhee]r}b  (h!]r~b  (h#h$e]rb  (h	j�  e]r�b  (hh�e]r�b  (h)h�eeejob  ]r�b  (j�^  ]r�b  (j�^  ]r�b  (j�^  ]r�b  (h	h�e]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	h�e]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	h
e]r�b  (hh<eeee]r�b  (hhee]r�b  (h!]r�b  (h#h$e]r�b  (h	j�  e]r�b  (hh�e]r�b  (h)h�eee]r�b  (j�^  ]r�b  (j�^  ]r�b  (j�^  ]r�b  (h	h�e]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	h�e]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	h
e]r�b  (hh<eeee]r�b  (hhee]r�b  (h!]r�b  (h#h$e]r�b  (h	j�  e]r�b  (hh�e]r�b  (h)h�eeej�b  ]r�b  (j�^  ]r�b  (j�^  ]r�b  (j�^  ]r�b  (h	h�e]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	h�e]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	h
e]r�b  (hh<eeee]r�b  (hhee]r�b  (h!]r�b  (h#h$e]r�b  (h	j�  e]r�b  (hh�e]r�b  (h)heee]r�b  (j�^  ]r�b  (j�^  ]r�b  (j�^  ]r�b  (h	h�e]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	he]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	h
e]r�b  (hh<eeee]r�b  (hhee]r�b  (h!]r�b  (h#h$e]r�b  (h	j�  e]r�b  (hh�e]r�b  (h)heee]r�b  (j�^  ]r�b  (j�^  ]r�b  (j�^  ]r�b  (h	h�e]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	he]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	h
e]r�b  (hh�eeee]r�b  (hhee]r�b  (h!]r�b  (h#h$e]r�b  (h	j�  e]r�b  (hh�e]r�b  (h)heee]r�b  (j�^  ]r�b  (j�^  ]r�b  (j�^  ]r�b  (h	h�e]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	he]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	h
e]r�b  (hh�eeee]r�b  (hhee]r�b  (h!]r�b  (h#h$e]r�b  (h	j�  e]r�b  (hh�e]r�b  (h)heeej�b  j�b  j�b  ]r�b  (j�^  ]r�b  (j�^  ]r�b  (j�^  ]r�b  (h	h�e]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	he]r�b  (hh�e]r�b  (hhe]r�b  (j�^  ]r�b  (h	h
e]r c  (hh�eeee]rc  (hhee]rc  (h!]rc  (h#h$e]rc  (h	j�  e]rc  (hh�e]rc  (h)heee]rc  (j�^  ]rc  (j�^  ]r	c  (j�^  ]r
c  (h	h�e]rc  (hh�e]rc  (hhe]rc  (j�^  ]rc  (h	he]rc  (hh�e]rc  (hhe]rc  (j�^  ]rc  (h	h
e]rc  (hh�eeee]rc  (hhee]rc  (h!]rc  (h#h$e]rc  (h	he]rc  (hh�e]rc  (h)h�eeejc  ]rc  (j�^  ]rc  (j�^  ]rc  (j�^  ]rc  (h	h�e]rc  (hh�e]rc  (hhe]r c  (j�^  ]r!c  (h	he]r"c  (hh�e]r#c  (hhe]r$c  (j�^  ]r%c  (h	h
e]r&c  (hh�eeee]r'c  (hhee]r(c  (h!]r)c  (h#h$e]r*c  (h	he]r+c  (hh�e]r,c  (h)h�eee]r-c  (j�^  ]r.c  (j�^  ]r/c  (j�^  ]r0c  (h	h�e]r1c  (hh�e]r2c  (hhe]r3c  (j�^  ]r4c  (h	he]r5c  (hh�e]r6c  (hhe]r7c  (j�^  ]r8c  (h	h
e]r9c  (hh�eeee]r:c  (hhee]r;c  (h!]r<c  (h#h$e]r=c  (h	he]r>c  (hh�e]r?c  (h)h�eeej-c  ]r@c  (j�^  ]rAc  (j�^  ]rBc  (j�^  ]rCc  (h	h�e]rDc  (hh�e]rEc  (hhe]rFc  (j�^  ]rGc  (h	he]rHc  (hh�e]rIc  (hhe]rJc  (j�^  ]rKc  (h	h
e]rLc  (hh�eeee]rMc  (hhee]rNc  (h!]rOc  (h#h$e]rPc  (h	he]rQc  (hh�e]rRc  (h)h�eeej@c  j@c  j@c  j@c  ]rSc  (j�^  ]rTc  (j�^  ]rUc  (j�^  ]rVc  (h	h�e]rWc  (hh�e]rXc  (hhe]rYc  (j�^  ]rZc  (h	he]r[c  (hh�e]r\c  (hhe]r]c  (j�^  ]r^c  (h	h�e]r_c  (hh�eeee]r`c  (hhee]rac  (h!]rbc  (h#h$e]rcc  (h	he]rdc  (hh�e]rec  (h)h�eeejSc  jSc  jSc  jSc  ]rfc  (j�^  ]rgc  (j�^  ]rhc  (j�^  ]ric  (h	h�e]rjc  (hh�e]rkc  (hhe]rlc  (j�^  ]rmc  (h	he]rnc  (hh�e]roc  (hhe]rpc  (j�^  ]rqc  (h	h�e]rrc  (hh�eeee]rsc  (hhee]rtc  (h!]ruc  (h#h$e]rvc  (h	he]rwc  (hh�e]rxc  (h)h�eeejfc  ]ryc  (j�^  ]rzc  (j�^  ]r{c  (j�^  ]r|c  (h	h�e]r}c  (hh�e]r~c  (hhe]rc  (j�^  ]r�c  (h	he]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�eeee]r�c  (hhee]r�c  (h!]r�c  (h#h$e]r�c  (h	he]r�c  (hh�e]r�c  (h)h�eee]r�c  (j�^  ]r�c  (j�^  ]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	he]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�eeee]r�c  (hhee]r�c  (h!]r�c  (h#h$e]r�c  (h	he]r�c  (hh�e]r�c  (h)h�eeej�c  ]r�c  (j�^  ]r�c  (j�^  ]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	he]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�eeee]r�c  (hhee]r�c  (h!]r�c  (h#h$e]r�c  (h	he]r�c  (hh�e]r�c  (h)h�eee]r�c  (j�^  ]r�c  (j�^  ]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	he]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�eeee]r�c  (hhee]r�c  (h!]r�c  (h#h$e]r�c  (h	he]r�c  (hh�e]r�c  (h)h�eeej�c  j�c  j�c  ]r�c  (j�^  ]r�c  (j�^  ]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	he]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�eeee]r�c  (hhee]r�c  (h!]r�c  (h#h$e]r�c  (h	he]r�c  (hh�e]r�c  (h)h�eeej�c  j�c  j�c  j�c  ]r�c  (j�^  ]r�c  (j�^  ]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	he]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�eeee]r�c  (hhee]r�c  (h!]r�c  (h#h$e]r�c  (h	he]r�c  (hh�e]r�c  (h)h�eee]r�c  (j�^  ]r�c  (j�^  ]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	he]r�c  (hh�e]r�c  (hhe]r�c  (j�^  ]r�c  (h	h�e]r�c  (hh�eeee]r�c  (hhee]r�c  (h!]r�c  (h#h$e]r�c  (h	he]r�c  (hh�e]r�c  (h)h�eeej�c  j�c  j�c  j�c  j�c  j�c  j�c  j�c  j�c  ]r�c  (j�^  ]r�c  (j�^  ]r d  (j�^  ]rd  (h	h�e]rd  (hh�e]rd  (hhe]rd  (j�^  ]rd  (h	he]rd  (hh�e]rd  (hhe]rd  (j�^  ]r	d  (h	h�e]r
d  (hh�eeee]rd  (hhee]rd  (h!]rd  (h#h$e]rd  (h	he]rd  (hh�e]rd  (h)h�eee]rd  (j�^  ]rd  (j�^  ]rd  (j�^  ]rd  (h	h�e]rd  (hh�e]rd  (hhe]rd  (j�^  ]rd  (h	he]rd  (hh�e]rd  (hhe]rd  (j�^  ]rd  (h	h�e]rd  (hh�eeee]rd  (hhee]rd  (h!]r d  (h#h$e]r!d  (h	he]r"d  (hh�e]r#d  (h)h�eeejd  jd  jd  ]r$d  (j�^  ]r%d  (j�^  ]r&d  (j�^  ]r'd  (h	h�e]r(d  (hh�e]r)d  (hhe]r*d  (j�^  ]r+d  (h	he]r,d  (hh�e]r-d  (hhe]r.d  (j�^  ]r/d  (h	h�e]r0d  (hh�eeee]r1d  (hhee]r2d  (h!]r3d  (h#h$e]r4d  (h	he]r5d  (hh�e]r6d  (h)h�eeej$d  ]r7d  (j�^  ]r8d  (j�^  ]r9d  (j�^  ]r:d  (h	h�e]r;d  (hh�e]r<d  (hhe]r=d  (j�^  ]r>d  (h	he]r?d  (hh�e]r@d  (hhe]rAd  (j�^  ]rBd  (h	h�e]rCd  (hh�eeee]rDd  (hhee]rEd  (h!]rFd  (h#h$e]rGd  (h	he]rHd  (hh�e]rId  (h)h�eeej7d  j7d  j7d  j7d  ]rJd  (j�^  ]rKd  (j�^  ]rLd  (j�^  ]rMd  (h	h�e]rNd  (hh�e]rOd  (hhe]rPd  (j�^  ]rQd  (h	he]rRd  (hh�e]rSd  (hhe]rTd  (j�^  ]rUd  (h	h�e]rVd  (hh�eeee]rWd  (hhee]rXd  (h!]rYd  (h#h$e]rZd  (h	he]r[d  (hh�e]r\d  (h)h�eee]r]d  (j�^  ]r^d  (j�^  ]r_d  (j�^  ]r`d  (h	h�e]rad  (hh�e]rbd  (hhe]rcd  (j�^  ]rdd  (h	he]red  (hh�e]rfd  (hhe]rgd  (j�^  ]rhd  (h	h�e]rid  (hh�eeee]rjd  (hhee]rkd  (h!]rld  (h#h$e]rmd  (h	he]rnd  (hh�e]rod  (h)h�eeej]d  ]rpd  (j�^  ]rqd  (j�^  ]rrd  (j�^  ]rsd  (h	h�e]rtd  (hh�e]rud  (hhe]rvd  (j�^  ]rwd  (h	he]rxd  (hh�e]ryd  (hhe]rzd  (j�^  ]r{d  (h	h�e]r|d  (hh�eeee]r}d  (hhee]r~d  (h!]rd  (h#h$e]r�d  (h	he]r�d  (hh�e]r�d  (h)h�eeejpd  jpd  jpd  jpd  jpd  jpd  jpd  jpd  jpd  jpd  jpd  jpd  jpd  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	he]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�eeee]r�d  (hhee]r�d  (h!]r�d  (h#h$e]r�d  (h	he]r�d  (hh�e]r�d  (h)h�eeej�d  j�d  j�d  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	he]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�eeee]r�d  (hhee]r�d  (h!]r�d  (h#h$e]r�d  (h	he]r�d  (hh�e]r�d  (h)h�eeej�d  j�d  j�d  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	he]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�eeee]r�d  (hhee]r�d  (h!]r�d  (h#h$e]r�d  (h	he]r�d  (hh�e]r�d  (h)h�eeej�d  j�d  j�d  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	he]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�eeee]r�d  (hhee]r�d  (h!]r�d  (h#h$e]r�d  (h	he]r�d  (hh�e]r�d  (h)h�eeej�d  j�d  j�d  j�d  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	he]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�eeee]r�d  (hhee]r�d  (h!]r�d  (h#h$e]r�d  (h	he]r�d  (hh�e]r�d  (h)h�eee]r�d  (j�^  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	he]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�eeee]r�d  (hhee]r�d  (h!]r�d  (h#h$e]r�d  (h	he]r�d  (hh�e]r�d  (h)h�eeej�d  j�d  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (j�^  ]r�d  (h	h�e]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r�d  (h	he]r�d  (hh�e]r�d  (hhe]r�d  (j�^  ]r e  (h	h�e]re  (hh�eeee]re  (hhee]re  (h!]re  (h#h$e]re  (h	he]re  (hh�e]re  (h)h�eeej�d  j�d  ]re  (j�^  ]r	e  (j�^  ]r
e  (j�^  ]re  (h	h�e]re  (hh�e]re  (hhe]re  (j�^  ]re  (h	he]re  (hh�e]re  (hhe]re  (j�^  ]re  (h	h�e]re  (hh�eeee]re  (hhee]re  (h!]re  (h#h$e]re  (h	he]re  (hh�e]re  (h)h�eee]re  (j�^  ]re  (j�^  ]re  (j�^  ]re  (h	h�e]re  (hh�e]r e  (hhe]r!e  (j�^  ]r"e  (h	he]r#e  (hh�e]r$e  (hhe]r%e  (j�^  ]r&e  (h	h�e]r'e  (hh�eeee]r(e  (hhee]r)e  (h!]r*e  (h#h$e]r+e  (h	he]r,e  (hh�e]r-e  (h)h�eee]r.e  (j�^  ]r/e  (j�^  ]r0e  (j�^  ]r1e  (h	h�e]r2e  (hh�e]r3e  (hhe]r4e  (j�^  ]r5e  (h	he]r6e  (hh�e]r7e  (hhe]r8e  (j�^  ]r9e  (h	h�e]r:e  (hh�eeee]r;e  (hhee]r<e  (h!]r=e  (h#h$e]r>e  (h	he]r?e  (hh�e]r@e  (h)h�eeej.e  j.e  j.e  j.e  j.e  ]rAe  (j�^  ]rBe  (j�^  ]rCe  (j�^  ]rDe  (h	h�e]rEe  (hh�e]rFe  (hhe]rGe  (j�^  ]rHe  (h	he]rIe  (hh�e]rJe  (hhe]rKe  (j�^  ]rLe  (h	h�e]rMe  (hh�eeee]rNe  (hhee]rOe  (h!]rPe  (h#h$e]rQe  (h	he]rRe  (hh�e]rSe  (h)h�eee]rTe  (j�^  ]rUe  (j�^  ]rVe  (j�^  ]rWe  (h	h�e]rXe  (hh�e]rYe  (hhe]rZe  (j�^  ]r[e  (h	he]r\e  (hh�e]r]e  (hhe]r^e  (j�^  ]r_e  (h	h�e]r`e  (hh�eeee]rae  (hhee]rbe  (h!]rce  (h#h$e]rde  (h	he]ree  (hh�e]rfe  (h)h�eeejTe  jTe  jTe  jTe  jTe  ]rge  (j�^  ]rhe  (j�^  ]rie  (j�^  ]rje  (h	h�e]rke  (hh�e]rle  (hhe]rme  (j�^  ]rne  (h	he]roe  (hh�e]rpe  (hhe]rqe  (j�^  ]rre  (h	h�e]rse  (hh�eeee]rte  (hhee]rue  (h!]rve  (h#h$e]rwe  (h	he]rxe  (hh�e]rye  (h)h�eee]rze  (j�^  ]r{e  (j�^  ]r|e  (j�^  ]r}e  (h	h�e]r~e  (hh�e]re  (hhe]r�e  (j�^  ]r�e  (h	he]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�eeee]r�e  (hhee]r�e  (h!]r�e  (h#h$e]r�e  (h	he]r�e  (hh�e]r�e  (h)h�eeejze  jze  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	he]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�eeee]r�e  (hhee]r�e  (h!]r�e  (h#h$e]r�e  (h	he]r�e  (hh�e]r�e  (h)h�eeej�e  j�e  j�e  j�e  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	he]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�eeee]r�e  (hhee]r�e  (h!]r�e  (h#h$e]r�e  (h	he]r�e  (hh�e]r�e  (h)h�eeej�e  j�e  j�e  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	he]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�eeee]r�e  (hhee]r�e  (h!]r�e  (h#h$e]r�e  (h	he]r�e  (hh�e]r�e  (h)h�eeej�e  j�e  j�e  j�e  j�e  j�e  j�e  j�e  j�e  j�e  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	he]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�eeee]r�e  (hhee]r�e  (h!]r�e  (h#h$e]r�e  (h	he]r�e  (hh�e]r�e  (h)h�eeej�e  j�e  j�e  j�e  j�e  j�e  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	he]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�eeee]r�e  (hhee]r�e  (h!]r�e  (h#h$e]r�e  (h	he]r�e  (hh�e]r�e  (h)h�eeej�e  j�e  j�e  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	he]r�e  (hh�e]r�e  (hhe]r�e  (j�^  ]r�e  (h	h�e]r�e  (hh�eeee]r�e  (hhee]r�e  (h!]r�e  (h#h$e]r�e  (h	he]r�e  (hh�e]r�e  (h)h�eeej�e  ]r�e  (j�^  ]r f  (j�^  ]rf  (j�^  ]rf  (h	h�e]rf  (hh�e]rf  (hhe]rf  (j�^  ]rf  (h	he]rf  (hh�e]rf  (hhe]r	f  (j�^  ]r
f  (h	h�e]rf  (hh�eeee]rf  (hhee]rf  (h!]rf  (h#h$e]rf  (h	he]rf  (hh�e]rf  (h)h�eeej�e  ]rf  (j�^  ]rf  (j�^  ]rf  (j�^  ]rf  (h	h�e]rf  (hh�e]rf  (hhe]rf  (j�^  ]rf  (h	he]rf  (hh�e]rf  (hhe]rf  (j�^  ]rf  (h	h�e]rf  (hh�eeee]rf  (hhee]r f  (h!]r!f  (h#h$e]r"f  (h	he]r#f  (hh�e]r$f  (h)h�eeejf  jf  ]r%f  (j�^  ]r&f  (j�^  ]r'f  (j�^  ]r(f  (h	h�e]r)f  (hh�e]r*f  (hhe]r+f  (j�^  ]r,f  (h	he]r-f  (hh�e]r.f  (hhe]r/f  (j�^  ]r0f  (h	h�e]r1f  (hh�eeee]r2f  (hhee]r3f  (h!]r4f  (h#h$e]r5f  (h	he]r6f  (hh�e]r7f  (h)h�eee]r8f  (j�^  ]r9f  (j�^  ]r:f  (j�^  ]r;f  (h	h�e]r<f  (hh�e]r=f  (hhe]r>f  (j�^  ]r?f  (h	he]r@f  (hh�e]rAf  (hhe]rBf  (j�^  ]rCf  (h	h�e]rDf  (hh�eeee]rEf  (hhee]rFf  (h!]rGf  (h#h$e]rHf  (h	he]rIf  (hh�e]rJf  (h)heeej8f  ]rKf  (j�^  ]rLf  (j�^  ]rMf  (j�^  ]rNf  (h	h�e]rOf  (hh�e]rPf  (hhe]rQf  (j�^  ]rRf  (h	he]rSf  (hh�e]rTf  (hhe]rUf  (j�^  ]rVf  (h	h�e]rWf  (hh�eeee]rXf  (hhee]rYf  (h!]rZf  (h#h$e]r[f  (h	he]r\f  (hh�e]r]f  (h)heeejKf  jKf  jKf  jKf  jKf  ]r^f  (j�^  ]r_f  (j�^  ]r`f  (j�^  ]raf  (h	h�e]rbf  (hh�e]rcf  (hhe]rdf  (j�^  ]ref  (h	he]rff  (hh�e]rgf  (hhe]rhf  (j�^  ]rif  (h	h�e]rjf  (hh�eeee]rkf  (hhee]rlf  (h!]rmf  (h#h$e]rnf  (h	he]rof  (hh�e]rpf  (h)heeej^f  j^f  ]rqf  (j�^  ]rrf  (j�^  ]rsf  (j�^  ]rtf  (h	h�e]ruf  (hh�e]rvf  (hhe]rwf  (j�^  ]rxf  (h	he]ryf  (hh�e]rzf  (hhe]r{f  (j�^  ]r|f  (h	h�e]r}f  (hh�eeee]r~f  (hhee]rf  (h!]r�f  (h#h$e]r�f  (h	he]r�f  (hh�e]r�f  (h)heeejqf  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	he]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�eeee]r�f  (hhee]r�f  (h!]r�f  (h#h$e]r�f  (h	he]r�f  (hh�e]r�f  (h)heee]r�f  (j�^  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	he]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�eeee]r�f  (hhee]r�f  (h!]r�f  (h#h$e]r�f  (h	he]r�f  (hh�e]r�f  (h)heeej�f  j�f  j�f  j�f  j�f  j�f  j�f  j�f  j�f  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	he]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�eeee]r�f  (hhee]r�f  (h!]r�f  (h#h$e]r�f  (h	he]r�f  (hh�e]r�f  (h)heeej�f  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	he]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�eeee]r�f  (hhee]r�f  (h!]r�f  (h#h$e]r�f  (h	he]r�f  (hh�e]r�f  (h)heeej�f  j�f  j�f  j�f  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	he]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�eeee]r�f  (hhee]r�f  (h!]r�f  (h#h$e]r�f  (h	he]r�f  (hh�e]r�f  (h)heeej�f  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	he]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�eeee]r�f  (hhee]r�f  (h!]r�f  (h#h$e]r�f  (h	he]r�f  (hh�e]r�f  (h)heee]r�f  (j�^  ]r�f  (j�^  ]r�f  (j�^  ]r�f  (h	h�e]r�f  (hh�e]r�f  (hhe]r�f  (j�^  ]r�f  (h	he]r�f  (hh�e]r�f  (hhe]r g  (j�^  ]rg  (h	h�e]rg  (hh�eeee]rg  (hhee]rg  (h!]rg  (h#h$e]rg  (h	he]rg  (hh�e]rg  (h)heeej�f  ]r	g  (j�^  ]r
g  (j�^  ]rg  (j�^  ]rg  (h	h�e]rg  (hh�e]rg  (hhe]rg  (j�^  ]rg  (h	he]rg  (hh�e]rg  (hhe]rg  (j�^  ]rg  (h	h�e]rg  (hh�eeee]rg  (hhee]rg  (h!]rg  (h#h$e]rg  (h	he]rg  (hh�e]rg  (h)heeej	g  j	g  j	g  j	g  j	g  j	g  j	g  j	g  j	g  ]rg  (j�^  ]rg  (j�^  ]rg  (j�^  ]rg  (h	h�e]r g  (hh�e]r!g  (hhe]r"g  (j�^  ]r#g  (h	he]r$g  (hh�e]r%g  (hhe]r&g  (j�^  ]r'g  (h	h�e]r(g  (hh�eeee]r)g  (hhee]r*g  (h!]r+g  (h#h$e]r,g  (h	he]r-g  (hh�e]r.g  (h)heeejg  jg  jg  ]r/g  (j�^  ]r0g  (j�^  ]r1g  (j�^  ]r2g  (h	h�e]r3g  (hh�e]r4g  (hhe]r5g  (j�^  ]r6g  (h	he]r7g  (hh�e]r8g  (hhe]r9g  (j�^  ]r:g  (h	h�e]r;g  (hh�eeee]r<g  (hhee]r=g  (h!]r>g  (h#h$e]r?g  (h	he]r@g  (hh�e]rAg  (h)heee]rBg  (j�^  ]rCg  (j�^  ]rDg  (j�^  ]rEg  (h	h�e]rFg  (hh�e]rGg  (hhe]rHg  (j�^  ]rIg  (h	he]rJg  (hh�e]rKg  (hhe]rLg  (j�^  ]rMg  (h	h�e]rNg  (hh�eeee]rOg  (hhee]rPg  (h!]rQg  (h#h$e]rRg  (h	he]rSg  (hh�e]rTg  (h)heee]rUg  (j�^  ]rVg  (j�^  ]rWg  (j�^  ]rXg  (h	h�e]rYg  (hh�e]rZg  (hhe]r[g  (j�^  ]r\g  (h	he]r]g  (hh�e]r^g  (hhe]r_g  (j�^  ]r`g  (h	h�e]rag  (hh�eeee]rbg  (hhee]rcg  (h!]rdg  (h#h$e]reg  (h	he]rfg  (hh�e]rgg  (h)heeejUg  ]rhg  (j�^  ]rig  (j�^  ]rjg  (j�^  ]rkg  (h	h�e]rlg  (hh�e]rmg  (hhe]rng  (j�^  ]rog  (h	he]rpg  (hh�e]rqg  (hhe]rrg  (j�^  ]rsg  (h	h�e]rtg  (hh�eeee]rug  (hhee]rvg  (h!]rwg  (h#h$e]rxg  (h	he]ryg  (hh�e]rzg  (h)heeejhg  ]r{g  (j�^  ]r|g  (j�^  ]r}g  (j�^  ]r~g  (h	h�e]rg  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	he]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�eeee]r�g  (hhee]r�g  (h!]r�g  (h#h$e]r�g  (h	he]r�g  (hh�e]r�g  (h)heeej{g  ]r�g  (j�^  ]r�g  (j�^  ]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	he]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�eeee]r�g  (hhee]r�g  (h!]r�g  (h#h$e]r�g  (h	he]r�g  (hh�e]r�g  (h)heee]r�g  (j�^  ]r�g  (j�^  ]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	he]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�eeee]r�g  (hhee]r�g  (h!]r�g  (h#h$e]r�g  (h	he]r�g  (hh�e]r�g  (h)heeej�g  ]r�g  (j�^  ]r�g  (j�^  ]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	he]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�eeee]r�g  (hhee]r�g  (h!]r�g  (h#h$e]r�g  (h	he]r�g  (hh�e]r�g  (h)heee]r�g  (j�^  ]r�g  (j�^  ]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	he]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�eeee]r�g  (hhee]r�g  (h!]r�g  (h#h$e]r�g  (h	he]r�g  (hh�e]r�g  (h)heeej�g  ]r�g  (j�^  ]r�g  (j�^  ]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	he]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�eeee]r�g  (hhee]r�g  (h!]r�g  (h#h$e]r�g  (h	he]r�g  (hh�e]r�g  (h)heee]r�g  (j�^  ]r�g  (j�^  ]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	he]r�g  (hh�e]r�g  (hhe]r�g  (j�^  ]r�g  (h	h�e]r�g  (hh�eeee]r�g  (hhee]r�g  (h!]r�g  (h#h$e]r�g  (h	he]r�g  (hh�e]r�g  (h)heee]r h  (j�^  ]rh  (j�^  ]rh  (j�^  ]rh  (h	h�e]rh  (hh�e]rh  (hhe]rh  (j�^  ]rh  (h	he]rh  (hh�e]r	h  (hhe]r
h  (j�^  ]rh  (h	h�e]rh  (hh�eeee]rh  (hhee]rh  (h!]rh  (h#h$e]rh  (h	he]rh  (hh�e]rh  (h)heee]rh  (j�^  ]rh  (j�^  ]rh  (j�^  ]rh  (h	h�e]rh  (hh�e]rh  (hhe]rh  (j�^  ]rh  (h	he]rh  (hh�e]rh  (hhe]rh  (j�^  ]rh  (h	h�e]rh  (hh�eeee]r h  (hhee]r!h  (h!]r"h  (h#h$e]r#h  (h	he]r$h  (hh�e]r%h  (h)heeejh  jh  jh  jh  jh  ]r&h  (j�^  ]r'h  (j�^  ]r(h  (j�^  ]r)h  (h	h�e]r*h  (hh�e]r+h  (hhe]r,h  (j�^  ]r-h  (h	he]r.h  (hh�e]r/h  (hhe]r0h  (j�^  ]r1h  (h	h�e]r2h  (hh�eeee]r3h  (hhee]r4h  (h!]r5h  (h#h$e]r6h  (h	he]r7h  (hh�e]r8h  (h)heeej&h  ]r9h  (j�^  ]r:h  (j�^  ]r;h  (j�^  ]r<h  (h	h�e]r=h  (hh�e]r>h  (hhe]r?h  (j�^  ]r@h  (h	he]rAh  (hh�e]rBh  (hhe]rCh  (j�^  ]rDh  (h	h�e]rEh  (hh�eeee]rFh  (hhee]rGh  (h!]rHh  (h#h$e]rIh  (h	he]rJh  (hh�e]rKh  (h)heeej9h  j9h  j9h  ]rLh  (j�^  ]rMh  (j�^  ]rNh  (j�^  ]rOh  (h	h�e]rPh  (hh�e]rQh  (hhe]rRh  (j�^  ]rSh  (h	he]rTh  (hh�e]rUh  (hhe]rVh  (j�^  ]rWh  (h	h�e]rXh  (hh�eeee]rYh  (hhee]rZh  (h!]r[h  (h#h$e]r\h  (h	he]r]h  (hh�e]r^h  (h)heeejLh  jLh  jLh  jLh  jLh  jLh  ]r_h  (j�^  ]r`h  (j�^  ]rah  (j�^  ]rbh  (h	h�e]rch  (hh�e]rdh  (hhe]reh  (j�^  ]rfh  (h	he]rgh  (hh�e]rhh  (hhe]rih  (j�^  ]rjh  (h	h�e]rkh  (hh�eeee]rlh  (hhee]rmh  (h!]rnh  (h#h$e]roh  (h	he]rph  (hh�e]rqh  (h)heeej_h  j_h  j_h  j_h  j_h  j_h  j_h  ]rrh  (j�^  ]rsh  (j�^  ]rth  (j�^  ]ruh  (h	h�e]rvh  (hh�e]rwh  (hhe]rxh  (j�^  ]ryh  (h	h�e]rzh  (hh�e]r{h  (hhe]r|h  (j�^  ]r}h  (h	h�e]r~h  (hh�eeee]rh  (hhee]r�h  (h!]r�h  (h#h$e]r�h  (h	he]r�h  (hh�e]r�h  (h)heeejrh  jrh  jrh  jrh  jrh  jrh  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�eeee]r�h  (hhee]r�h  (h!]r�h  (h#h$e]r�h  (h	he]r�h  (hh�e]r�h  (h)heeej�h  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�eeee]r�h  (hhee]r�h  (h!]r�h  (h#h$e]r�h  (h	he]r�h  (hh�e]r�h  (h)heeej�h  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�eeee]r�h  (hhee]r�h  (h!]r�h  (h#h$e]r�h  (h	he]r�h  (hh�e]r�h  (h)heeej�h  j�h  j�h  j�h  j�h  j�h  j�h  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�eeee]r�h  (hhee]r�h  (h!]r�h  (h#h$e]r�h  (h	he]r�h  (hh�e]r�h  (h)heeej�h  j�h  j�h  j�h  j�h  j�h  j�h  j�h  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�eeee]r�h  (hhee]r�h  (h!]r�h  (h#h$e]r�h  (h	he]r�h  (hh�e]r�h  (h)heee]r�h  (j�^  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�eeee]r�h  (hhee]r�h  (h!]r�h  (h#h$e]r�h  (h	he]r�h  (hh�e]r�h  (h)heeej�h  j�h  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r�h  (hhe]r�h  (j�^  ]r�h  (h	h�e]r�h  (hh�e]r i  (hhe]ri  (j�^  ]ri  (h	h�e]ri  (hh�eeee]ri  (hhee]ri  (h!]ri  (h#h$e]ri  (h	he]ri  (hh�e]r	i  (h)heee]r
i  (j�^  ]ri  (j�^  ]ri  (j�^  ]ri  (h	h�e]ri  (hh�e]ri  (hhe]ri  (j�^  ]ri  (h	h�e]ri  (hh�e]ri  (hhe]ri  (j�^  ]ri  (h	h�e]ri  (hh�eeee]ri  (hhee]ri  (h!]ri  (h#h$e]ri  (h	he]ri  (hh�e]ri  (h)heee]ri  (j�^  ]ri  (j�^  ]ri  (j�^  ]r i  (h	h�e]r!i  (hh�e]r"i  (hhe]r#i  (j�^  ]r$i  (h	h�e]r%i  (hh�e]r&i  (hhe]r'i  (j�^  ]r(i  (h	h�e]r)i  (hh�eeee]r*i  (hhee]r+i  (h!]r,i  (h#h$e]r-i  (h	he]r.i  (hh�e]r/i  (h)heeeji  ji  ji  ]r0i  (j�^  ]r1i  (j�^  ]r2i  (j�^  ]r3i  (h	h�e]r4i  (hh�e]r5i  (hhe]r6i  (j�^  ]r7i  (h	h�e]r8i  (hh�e]r9i  (hhe]r:i  (j�^  ]r;i  (h	h�e]r<i  (hh�eeee]r=i  (hhee]r>i  (h!]r?i  (h#h$e]r@i  (h	he]rAi  (hh�e]rBi  (h)heeej0i  ]rCi  (j�^  ]rDi  (j�^  ]rEi  (j�^  ]rFi  (h	h�e]rGi  (hh�e]rHi  (hhe]rIi  (j�^  ]rJi  (h	h�e]rKi  (hh�e]rLi  (hhe]rMi  (j�^  ]rNi  (h	h�e]rOi  (hh�eeee]rPi  (hhee]rQi  (h!]rRi  (h#h$e]rSi  (h	he]rTi  (hh�e]rUi  (h)heee]rVi  (j�^  ]rWi  (j�^  ]rXi  (j�^  ]rYi  (h	h�e]rZi  (hh�e]r[i  (hhe]r\i  (j�^  ]r]i  (h	h�e]r^i  (hh�e]r_i  (hhe]r`i  (j�^  ]rai  (h	h�e]rbi  (hh�eeee]rci  (hhee]rdi  (h!]rei  (h#h$e]rfi  (h	he]rgi  (hh�e]rhi  (h)heeejVi  jVi  jVi  ]rii  (j�^  ]rji  (j�^  ]rki  (j�^  ]rli  (h	h�e]rmi  (hh�e]rni  (hhe]roi  (j�^  ]rpi  (h	h�e]rqi  (hh�e]rri  (hhe]rsi  (j�^  ]rti  (h	h�e]rui  (hh�eeee]rvi  (hhee]rwi  (h!]rxi  (h#h$e]ryi  (h	he]rzi  (hh�e]r{i  (h)heeejii  jii  jii  jii  ]r|i  (j�^  ]r}i  (j�^  ]r~i  (j�^  ]ri  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�eeee]r�i  (hhee]r�i  (h!]r�i  (h#h$e]r�i  (h	he]r�i  (hh�e]r�i  (h)heeej|i  j|i  ]r�i  (j�^  ]r�i  (j�^  ]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�eeee]r�i  (hhee]r�i  (h!]r�i  (h#h$e]r�i  (h	he]r�i  (hh�e]r�i  (h)heee]r�i  (j�^  ]r�i  (j�^  ]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�eeee]r�i  (hhee]r�i  (h!]r�i  (h#h$e]r�i  (h	he]r�i  (hh�e]r�i  (h)heeej�i  ]r�i  (j�^  ]r�i  (j�^  ]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�eeee]r�i  (hhee]r�i  (h!]r�i  (h#h$e]r�i  (h	he]r�i  (hh�e]r�i  (h)heee]r�i  (j�^  ]r�i  (j�^  ]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (X	   Next-Mover�i  ]r�i  (h	h�e]r�i  (hh�eeee]r�i  (hhee]r�i  (h!]r�i  (h#h$e]r�i  (h	he]r�i  (hh�e]r�i  (h)heee]r�i  (j�^  ]r�i  (j�^  ]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�i  ]r�i  (h	h�e]r�i  (hh�eeee]r�i  (hhee]r�i  (h!]r�i  (h#h$e]r�i  (h	he]r�i  (hh�e]r�i  (h)heeej�i  j�i  j�i  ]r�i  (j�^  ]r�i  (j�^  ]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�^  ]r�i  (h	h�e]r�i  (hh�e]r�i  (hhe]r�i  (j�i  ]r�i  (h	h�e]r�i  (hh�eeee]r�i  (hhee]r�i  (h!]r�i  (h#h$e]r�i  (h	he]r j  (hh�e]rj  (h)heeej�i  j�i  j�i  j�i  j�i  j�i  j�i  j�i  j�i  j�i  j�i  j�i  j�i  ]rj  (j�^  ]rj  (j�^  ]rj  (j�^  ]rj  (h	h�e]rj  (hh�e]rj  (hhe]rj  (j�^  ]r	j  (h	h�e]r
j  (hh�e]rj  (hhe]rj  (j�i  ]rj  (h	h�e]rj  (hh�eeee]rj  (hhee]rj  (h!]rj  (h#h$e]rj  (h	he]rj  (hh�e]rj  (h)heeejj  jj  ]rj  (j�^  ]rj  (j�^  ]rj  (j�^  ]rj  (h	h�e]rj  (hh�e]rj  (hhe]rj  (j�^  ]rj  (h	he]rj  (hh�e]rj  (hhe]rj  (j�i  ]r j  (h	h�e]r!j  (hh�eeee]r"j  (hhee]r#j  (h!]r$j  (h#h$e]r%j  (h	he]r&j  (hh�e]r'j  (h)heeejj  jj  jj  ]r(j  (j�^  ]r)j  (j�^  ]r*j  (j�^  ]r+j  (h	h�e]r,j  (hh�e]r-j  (hhe]r.j  (j�^  ]r/j  (h	he]r0j  (hh�e]r1j  (hhe]r2j  (j�i  ]r3j  (h	h�e]r4j  (hh�eeee]r5j  (hhee]r6j  (h!]r7j  (h#h$e]r8j  (h	he]r9j  (hh�e]r:j  (h)heee]r;j  (j�^  ]r<j  (j�^  ]r=j  (j�^  ]r>j  (h	h�e]r?j  (hh�e]r@j  (hhe]rAj  (j�^  ]rBj  (h	he]rCj  (hh�e]rDj  (hhe]rEj  (j�i  ]rFj  (h	h�e]rGj  (hh�eeee]rHj  (hhee]rIj  (h!]rJj  (h#h$e]rKj  (h	he]rLj  (hh�e]rMj  (h)heee]rNj  (j�^  ]rOj  (j�^  ]rPj  (j�^  ]rQj  (h	h�e]rRj  (hh�e]rSj  (hhe]rTj  (j�^  ]rUj  (h	he]rVj  (hh�e]rWj  (hhe]rXj  (j�i  ]rYj  (h	h�e]rZj  (hh�eeee]r[j  (hhee]r\j  (h!]r]j  (h#h$e]r^j  (h	he]r_j  (hh�e]r`j  (h)heeejNj  jNj  ]raj  (j�^  ]rbj  (j�^  ]rcj  (j�^  ]rdj  (h	h�e]rej  (hh�e]rfj  (hhe]rgj  (j�^  ]rhj  (h	he]rij  (hh�e]rjj  (hhe]rkj  (j�i  ]rlj  (h	h�e]rmj  (hh�eeee]rnj  (hhee]roj  (h!]rpj  (h#h$e]rqj  (h	he]rrj  (hh�e]rsj  (h)heeejaj  jaj  jaj  jaj  jaj  jaj  jaj  jaj  jaj  jaj  jaj  jaj  jaj  jaj  jaj  jaj  ]rtj  (j�^  ]ruj  (j�^  ]rvj  (j�^  ]rwj  (h	h�e]rxj  (hh�e]ryj  (hhe]rzj  (j�^  ]r{j  (h	he]r|j  (hh�e]r}j  (hhe]r~j  (j�i  ]rj  (h	h�e]r�j  (hh�eeee]r�j  (hhee]r�j  (h!]r�j  (h#h$e]r�j  (h	he]r�j  (hh�e]r�j  (h)heeejtj  jtj  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (h	h�e]r�j  (hh�e]r�j  (hhe]r�j  (j�^  ]r�j  (h	he]r�j  (hh�e]r�j  (hhe]r�j  (j�i  ]r�j  (h	h�e]r�j  (hh�eeee]r�j  (hhee]r�j  (h!]r�j  (h#h$e]r�j  (h	he]r�j  (hh�e]r�j  (h)heee]r�j  (j�^  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (h	h�e]r�j  (hh�e]r�j  (hhe]r�j  (j�^  ]r�j  (h	he]r�j  (hh�e]r�j  (hhe]r�j  (j�i  ]r�j  (h	h�e]r�j  (hh�eeee]r�j  (hhee]r�j  (h!]r�j  (h#h$e]r�j  (h	he]r�j  (hh�e]r�j  (h)heee]r�j  (j�^  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (h	h�e]r�j  (hh�e]r�j  (hhe]r�j  (j�^  ]r�j  (h	he]r�j  (hh�e]r�j  (hhe]r�j  (j�i  ]r�j  (h	h�e]r�j  (hh�eeee]r�j  (hhee]r�j  (h!]r�j  (h#h$e]r�j  (h	he]r�j  (hh�e]r�j  (h)heeej�j  j�j  j�j  j�j  j�j  j�j  j�j  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (h	h�e]r�j  (hh�e]r�j  (hhe]r�j  (j�^  ]r�j  (h	he]r�j  (hh�e]r�j  (hhe]r�j  (j�i  ]r�j  (h	h�e]r�j  (hh�eeee]r�j  (hhee]r�j  (h!]r�j  (h#h$e]r�j  (h	he]r�j  (hh�e]r�j  (h)heeej�j  j�j  j�j  j�j  j�j  j�j  j�j  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (h	h�e]r�j  (hh�e]r�j  (hhe]r�j  (j�^  ]r�j  (h	he]r�j  (hh�e]r�j  (hhe]r�j  (j�i  ]r�j  (h	h�e]r�j  (hh�eeee]r�j  (hhee]r�j  (h!]r�j  (h#h$e]r�j  (h	he]r�j  (hh�e]r�j  (h)heeej�j  j�j  j�j  j�j  j�j  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (h	h�e]r�j  (hh�e]r�j  (hhe]r�j  (j�^  ]r�j  (h	he]r�j  (hh�e]r�j  (hhe]r�j  (j�i  ]r�j  (h	h�e]r�j  (hh�eeee]r�j  (hhee]r�j  (h!]r�j  (h#h$e]r�j  (h	he]r�j  (hh�e]r�j  (h)heeej�j  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (j�^  ]r�j  (h	h�e]r�j  (hh�e]r�j  (hhe]r�j  (j�^  ]r k  (h	he]rk  (hh�e]rk  (hhe]rk  (j�i  ]rk  (h	h�e]rk  (hh�eeee]rk  (hhee]rk  (h!]rk  (h#h$e]r	k  (h	he]r
k  (hh�e]rk  (h)heeej�j  ]rk  (j�^  ]rk  (j�^  ]rk  (j�^  ]rk  (h	h�e]rk  (hh�e]rk  (hhe]rk  (j�^  ]rk  (h	h�e]rk  (hh�e]rk  (hhe]rk  (j�i  ]rk  (h	h�e]rk  (hh�eeee]rk  (hhee]rk  (h!]rk  (h#h$e]rk  (h	he]rk  (hh�e]rk  (h)heeejk  jk  jk  jk  jk  ]rk  (j�^  ]r k  (j�^  ]r!k  (j�^  ]r"k  (h	h�e]r#k  (hh�e]r$k  (hhe]r%k  (j�^  ]r&k  (h	h�e]r'k  (hh�e]r(k  (hhe]r)k  (j�i  ]r*k  (h	h�e]r+k  (hh�eeee]r,k  (hhee]r-k  (h!]r.k  (h#h$e]r/k  (h	he]r0k  (hh�e]r1k  (h)heee]r2k  (j�^  ]r3k  (j�^  ]r4k  (j�^  ]r5k  (h	h�e]r6k  (hh�e]r7k  (hhe]r8k  (j�^  ]r9k  (h	h�e]r:k  (hh�e]r;k  (hhe]r<k  (j�i  ]r=k  (h	h�e]r>k  (hh�eeee]r?k  (hhee]r@k  (h!]rAk  (h#h$e]rBk  (h	he]rCk  (hh�e]rDk  (h)heeej2k  j2k  j2k  j2k  j2k  j2k  j2k  j2k  j2k  j2k  ]rEk  (j�^  ]rFk  (j�^  ]rGk  (j�^  ]rHk  (h	h�e]rIk  (hh�e]rJk  (hhe]rKk  (j�^  ]rLk  (h	he]rMk  (hh�e]rNk  (hhe]rOk  (j�i  ]rPk  (h	h�e]rQk  (hh�eeee]rRk  (hhee]rSk  (h!]rTk  (h#h$e]rUk  (h	he]rVk  (hh�e]rWk  (h)heeejEk  ]rXk  (j�^  ]rYk  (j�^  ]rZk  (j�^  ]r[k  (h	h�e]r\k  (hh�e]r]k  (hhe]r^k  (j�^  ]r_k  (h	he]r`k  (hh�e]rak  (hhe]rbk  (j�i  ]rck  (h	h�e]rdk  (hh�eeee]rek  (hhee]rfk  (h!]rgk  (h#h$e]rhk  (h	he]rik  (hh�e]rjk  (h)heee]rkk  (j�^  ]rlk  (j�^  ]rmk  (j�^  ]rnk  (h	h�e]rok  (hh�e]rpk  (hhe]rqk  (j�^  ]rrk  (h	he]rsk  (hh�e]rtk  (hhe]ruk  (j�i  ]rvk  (h	h�e]rwk  (hh�eeee]rxk  (hhee]ryk  (h!]rzk  (h#h$e]r{k  (h	he]r|k  (hh�e]r}k  (h)heeejkk  jkk  jkk  ]r~k  (j�^  ]rk  (j�^  ]r�k  (j�^  ]r�k  (h	h�e]r�k  (hh�e]r�k  (hhe]r�k  (j�^  ]r�k  (h	he]r�k  (hh�e]r�k  (hhe]r�k  (j�i  ]r�k  (h	h�e]r�k  (hh�eeee]r�k  (hhee]r�k  (h!]r�k  (h#h$e]r�k  (h	he]r�k  (hh�e]r�k  (h)heeej~k  j~k  j~k  j~k  j~k  j~k  ]r�k  (j�^  ]r�k  (j�^  ]r�k  (j�^  ]r�k  (h	h�e]r�k  (hh�e]r�k  (hhe]r�k  (j�^  ]r�k  (h	he]r�k  (hh�e]r�k  (hhe]r�k  (j�i  ]r�k  (h	h�e]r�k  (hh�eeee]r�k  (hhee]r�k  (h!]r�k  (h#h$e]r�k  (h	he]r�k  (hh�e]r�k  (h)heeej�k  j�k  ]r�k  (j�^  ]r�k  (j�^  ]r�k  (j�^  ]r�k  (h	h�e]r�k  (hh�e]r�k  (hhe]r�k  (j�^  ]r�k  (h	he]r�k  (hh�e]r�k  (hhe]r�k  (j�i  ]r�k  (h	h�e]r�k  (hh�eeee]r�k  (hhee]r�k  (h!]r�k  (h#h$e]r�k  (h	he]r�k  (hh�e]r�k  (h)heee]r�k  (j�^  ]r�k  (j�^  ]r�k  (j�^  ]r�k  (h	h�e]r�k  (hh�e]r�k  (hhe]r�k  (j�^  ]r�k  (h	he]r�k  (hh�e]r�k  (hhe]r�k  (j�i  ]r�k  (h	h�e]r�k  (hh�eeee]r�k  (hhee]r�k  (h!]r�k  (h#h$e]r�k  (h	he]r�k  (hh�e]r�k  (h)heeej�k  j�k  ]r�k  (j�^  ]r�k  (j�^  ]r�k  (j�^  ]r�k  (h	h�e]r�k  (hh�e]r�k  (hhe]r�k  (j�^  ]r�k  (h	he]r�k  (hh�e]r�k  (hhe]r�k  (j�i  ]r�k  (h	h�e]r�k  (hh�eeee]r�k  (hhee]r�k  (h!]r�k  (h#h$e]r�k  (h	he]r�k  (hh�e]r�k  (h)heeej�k  j�k  ]r�k  (j�^  ]r�k  (j�^  ]r�k  (j�^  ]r�k  (h	h�e]r�k  (hh�e]r�k  (hhe]r�k  (j�^  ]r�k  (h	he]r�k  (hh�e]r�k  (hhe]r�k  (j�i  ]r�k  (h	h�e]r�k  (hh�eeee]r�k  (hhee]r�k  (h!]r�k  (h#h$e]r�k  (h	he]r�k  (hh�e]r�k  (h)heeej�k  ]r�k  (j�^  ]r�k  (j�^  ]r�k  (j�^  ]r�k  (h	h�e]r�k  (hh�e]r�k  (hhe]r�k  (j�^  ]r�k  (h	he]r�k  (hh�e]r�k  (hhe]r�k  (j�i  ]r�k  (h	h�e]r�k  (hh�eeee]r�k  (hhee]r�k  (h!]r�k  (h#h$e]r l  (h	he]rl  (hh�e]rl  (h)heee]rl  (j�^  ]rl  (j�^  ]rl  (j�^  ]rl  (h	h�e]rl  (hh�e]rl  (hhe]r	l  (j�^  ]r
l  (h	he]rl  (hh�e]rl  (hhe]rl  (j�i  ]rl  (h	h�e]rl  (hh�eeee]rl  (hhee]rl  (h!]rl  (h#h$e]rl  (h	he]rl  (hh�e]rl  (h)heeejl  jl  jl  jl  ]rl  (j�^  ]rl  (j�^  ]rl  (j�^  ]rl  (h	h�e]rl  (hh�e]rl  (hhe]rl  (j�^  ]rl  (h	he]rl  (hh�e]rl  (hhe]r l  (j�i  ]r!l  (h	h�e]r"l  (hh�eeee]r#l  (hhee]r$l  (h!]r%l  (h#h$e]r&l  (h	he]r'l  (hh�e]r(l  (h)heeejl  jl  ]r)l  (j�^  ]r*l  (j�^  ]r+l  (j�^  ]r,l  (h	h�e]r-l  (hh�e]r.l  (hhe]r/l  (j�^  ]r0l  (h	he]r1l  (hh�e]r2l  (hhe]r3l  (j�i  ]r4l  (h	h�e]r5l  (hh�eeee]r6l  (hhee]r7l  (h!]r8l  (h#h$e]r9l  (h	he]r:l  (hh�e]r;l  (h)heeej)l  j)l  j)l  ]r<l  (j�^  ]r=l  (j�^  ]r>l  (j�^  ]r?l  (h	h�e]r@l  (hh�e]rAl  (hhe]rBl  (j�^  ]rCl  (h	h�e]rDl  (hh�e]rEl  (hhe]rFl  (j�i  ]rGl  (h	h�e]rHl  (hh�eeee]rIl  (hhee]rJl  (h!]rKl  (h#h$e]rLl  (h	he]rMl  (hh�e]rNl  (h)heeej<l  ]rOl  (j�^  ]rPl  (j�^  ]rQl  (j�^  ]rRl  (h	h�e]rSl  (hh�e]rTl  (hhe]rUl  (j�^  ]rVl  (h	h�e]rWl  (hh�e]rXl  (hhe]rYl  (j�i  ]rZl  (h	h�e]r[l  (hh�eeee]r\l  (hhee]r]l  (h!]r^l  (h#h$e]r_l  (h	he]r`l  (hh�e]ral  (h)heeejOl  jOl  jOl  jOl  ]rbl  (j�^  ]rcl  (j�^  ]rdl  (j�^  ]rel  (h	h�e]rfl  (hh�e]rgl  (hhe]rhl  (j�^  ]ril  (h	h�e]rjl  (hh�e]rkl  (hhe]rll  (j�i  ]rml  (h	h�e]rnl  (hh�eeee]rol  (hhee]rpl  (h!]rql  (h#h$e]rrl  (h	he]rsl  (hh�e]rtl  (h)heeejbl  jbl  jbl  ]rul  (j�^  ]rvl  (j�^  ]rwl  (j�^  ]rxl  (h	h�e]ryl  (hh�e]rzl  (hhe]r{l  (j�^  ]r|l  (h	h�e]r}l  (hh�e]r~l  (hhe]rl  (j�i  ]r�l  (h	h�e]r�l  (hh�eeee]r�l  (hhee]r�l  (h!]r�l  (h#h$e]r�l  (h	he]r�l  (hh�e]r�l  (h)heee]r�l  (j�^  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�i  ]r�l  (h	h�e]r�l  (hh�eeee]r�l  (hhee]r�l  (h!]r�l  (h#h$e]r�l  (h	he]r�l  (hh�e]r�l  (h)heeej�l  j�l  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�i  ]r�l  (h	h�e]r�l  (hh�eeee]r�l  (hhee]r�l  (h!]r�l  (h#h$e]r�l  (h	he]r�l  (hh�e]r�l  (h)heee]r�l  (j�^  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�i  ]r�l  (h	h�e]r�l  (hh�eeee]r�l  (hhee]r�l  (h!]r�l  (h#h$e]r�l  (h	he]r�l  (hh�e]r�l  (h)heeej�l  j�l  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�i  ]r�l  (h	h�e]r�l  (hh�eeee]r�l  (hhee]r�l  (h!]r�l  (h#h$e]r�l  (h	he]r�l  (hh�e]r�l  (h)heeej�l  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�i  ]r�l  (h	h�e]r�l  (hh�eeee]r�l  (hhee]r�l  (h!]r�l  (h#h$e]r�l  (h	he]r�l  (hh�e]r�l  (h)heeej�l  j�l  j�l  j�l  j�l  j�l  j�l  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r�l  (j�i  ]r�l  (h	h�e]r�l  (hh�eeee]r�l  (hhee]r�l  (h!]r�l  (h#h$e]r�l  (h	he]r�l  (hh�e]r�l  (h)heeej�l  j�l  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (j�^  ]r�l  (h	h�e]r�l  (hh�e]r�l  (hhe]r m  (j�^  ]rm  (h	h�e]rm  (hh�e]rm  (hhe]rm  (j�i  ]rm  (h	h�e]rm  (hh�eeee]rm  (hhee]rm  (h!]r	m  (h#h$e]r
m  (h	he]rm  (hh�e]rm  (h)heeej�l  j�l  j�l  ]rm  (j�^  ]rm  (j�^  ]rm  (j�^  ]rm  (h	h�e]rm  (hh�e]rm  (hhe]rm  (j�^  ]rm  (h	h�e]rm  (hh�e]rm  (hhe]rm  (j�i  ]rm  (h	h�e]rm  (hh�eeee]rm  (hhee]rm  (h!]rm  (h#h$e]rm  (h	he]rm  (hh�e]rm  (h)heeejm  jm  jm  jm  jm  jm  ]r m  (j�^  ]r!m  (j�^  ]r"m  (j�^  ]r#m  (h	h�e]r$m  (hh�e]r%m  (hhe]r&m  (j�^  ]r'm  (h	h�e]r(m  (hh�e]r)m  (hhe]r*m  (j�i  ]r+m  (h	h�e]r,m  (hh�eeee]r-m  (hhee]r.m  (h!]r/m  (h#h$e]r0m  (h	he]r1m  (hh�e]r2m  (h)heee]r3m  (j�^  ]r4m  (j�^  ]r5m  (j�^  ]r6m  (h	h�e]r7m  (hh�e]r8m  (hhe]r9m  (j�^  ]r:m  (h	h�e]r;m  (hh�e]r<m  (hhe]r=m  (j�i  ]r>m  (h	h�e]r?m  (hh�eeee]r@m  (hhee]rAm  (h!]rBm  (h#h$e]rCm  (h	he]rDm  (hh�e]rEm  (h)heeej3m  j3m  j3m  ]rFm  (j�^  ]rGm  (j�^  ]rHm  (j�^  ]rIm  (h	h�e]rJm  (hh�e]rKm  (hhe]rLm  (j�^  ]rMm  (h	h�e]rNm  (hh�e]rOm  (hhe]rPm  (j�i  ]rQm  (h	h�e]rRm  (hh�eeee]rSm  (hhee]rTm  (h!]rUm  (h#h$e]rVm  (h	he]rWm  (hh�e]rXm  (h)heeejFm  jFm  ]rYm  (j�^  ]rZm  (j�^  ]r[m  (j�^  ]r\m  (h	h�e]r]m  (hh�e]r^m  (hhe]r_m  (j�^  ]r`m  (h	h�e]ram  (hh�e]rbm  (hhe]rcm  (j�i  ]rdm  (h	h�e]rem  (hh�eeee]rfm  (hhee]rgm  (h!]rhm  (h#h$e]rim  (h	he]rjm  (hh�e]rkm  (h)heeejYm  jYm  ]rlm  (j�^  ]rmm  (j�^  ]rnm  (j�^  ]rom  (h	h�e]rpm  (hh�e]rqm  (hhe]rrm  (j�^  ]rsm  (h	h�e]rtm  (hh�e]rum  (hhe]rvm  (j�i  ]rwm  (h	h�e]rxm  (hh�eeee]rym  (hhee]rzm  (h!]r{m  (h#h$e]r|m  (h	he]r}m  (hh�e]r~m  (h)heeejlm  jlm  jlm  jlm  jlm  jlm  ]rm  (j�^  ]r�m  (j�^  ]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�i  ]r�m  (h	h�e]r�m  (hh�eeee]r�m  (hhee]r�m  (h!]r�m  (h#h$e]r�m  (h	he]r�m  (hh�e]r�m  (h)heee]r�m  (j�^  ]r�m  (j�^  ]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�i  ]r�m  (h	h�e]r�m  (hh�eeee]r�m  (hhee]r�m  (h!]r�m  (h#h$e]r�m  (h	he]r�m  (hh�e]r�m  (h)heeej�m  ]r�m  (j�^  ]r�m  (j�^  ]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�i  ]r�m  (h	h�e]r�m  (hh�eeee]r�m  (hhee]r�m  (h!]r�m  (h#h$e]r�m  (h	he]r�m  (hh�e]r�m  (h)heee]r�m  (j�^  ]r�m  (j�^  ]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�i  ]r�m  (h	h�e]r�m  (hh�eeee]r�m  (hhee]r�m  (h!]r�m  (h#h$e]r�m  (h	he]r�m  (hh�e]r�m  (h)heeej�m  j�m  j�m  j�m  j�m  ]r�m  (j�^  ]r�m  (j�^  ]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�i  ]r�m  (h	h�e]r�m  (hh�eeee]r�m  (hhee]r�m  (h!]r�m  (h#h$e]r�m  (h	he]r�m  (hh�e]r�m  (h)heee]r�m  (j�^  ]r�m  (j�^  ]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�^  ]r�m  (h	he]r�m  (hh�e]r�m  (hhe]r�m  (j�i  ]r�m  (h	h�e]r�m  (hh�eeee]r�m  (hhee]r�m  (h!]r�m  (h#h$e]r�m  (h	he]r�m  (hh�e]r�m  (h)heeej�m  j�m  ]r�m  (j�^  ]r�m  (j�^  ]r�m  (j�^  ]r�m  (h	h�e]r�m  (hh�e]r�m  (hhe]r�m  (j�^  ]r�m  (h	he]r�m  (hh�e]r�m  (hhe]r�m  (j�i  ]r�m  (h	h�e]r�m  (hh�eeee]r�m  (hhee]r�m  (h!]r n  (h#h$e]rn  (h	he]rn  (hh�e]rn  (h)heee]rn  (j�^  ]rn  (j�^  ]rn  (j�^  ]rn  (h	h�e]rn  (hh�e]r	n  (hhe]r
n  (j�^  ]rn  (h	he]rn  (hh�e]rn  (hhe]rn  (j�i  ]rn  (h	h�e]rn  (hh�eeee]rn  (hhee]rn  (h!]rn  (h#h$e]rn  (h	he]rn  (hh�e]rn  (h)heee]rn  (j�^  ]rn  (j�^  ]rn  (j�^  ]rn  (h	h�e]rn  (hh�e]rn  (hhe]rn  (j�^  ]rn  (h	he]rn  (hh�e]r n  (hhe]r!n  (j�i  ]r"n  (h	h�e]r#n  (hh�eeee]r$n  (hhee]r%n  (h!]r&n  (h#h$e]r'n  (h	he]r(n  (hh�e]r)n  (h)heeejn  ]r*n  (j�^  ]r+n  (j�^  ]r,n  (j�^  ]r-n  (h	h�e]r.n  (hh�e]r/n  (hhe]r0n  (j�^  ]r1n  (h	he]r2n  (hh�e]r3n  (hhe]r4n  (j�i  ]r5n  (h	h�e]r6n  (hh�eeee]r7n  (hhee]r8n  (h!]r9n  (h#h$e]r:n  (h	he]r;n  (hh�e]r<n  (h)heeej*n  j*n  j*n  j*n  j*n  j*n  ]r=n  (j�^  ]r>n  (j�^  ]r?n  (j�^  ]r@n  (h	h�e]rAn  (hh�e]rBn  (hhe]rCn  (j�^  ]rDn  (h	he]rEn  (hh�e]rFn  (hhe]rGn  (j�i  ]rHn  (h	h�e]rIn  (hh�eeee]rJn  (hhee]rKn  (h!]rLn  (h#h$e]rMn  (h	he]rNn  (hh�e]rOn  (h)heeej=n  ]rPn  (j�^  ]rQn  (j�^  ]rRn  (j�^  ]rSn  (h	h�e]rTn  (hh�e]rUn  (hhe]rVn  (j�^  ]rWn  (h	he]rXn  (hh�e]rYn  (hhe]rZn  (j�i  ]r[n  (h	h�e]r\n  (hh�eeee]r]n  (hhee]r^n  (h!]r_n  (h#h$e]r`n  (h	he]ran  (hh�e]rbn  (h)heeejPn  ]rcn  (j�^  ]rdn  (j�^  ]ren  (j�^  ]rfn  (h	h�e]rgn  (hh�e]rhn  (hhe]rin  (j�^  ]rjn  (h	he]rkn  (hh�e]rln  (hhe]rmn  (j�i  ]rnn  (h	h�e]ron  (hh�eeee]rpn  (hhee]rqn  (h!]rrn  (h#h$e]rsn  (h	he]rtn  (hh�e]run  (h)heeejcn  jcn  jcn  jcn  jcn  ]rvn  (j�^  ]rwn  (j�^  ]rxn  (j�^  ]ryn  (h	h�e]rzn  (hh�e]r{n  (hhe]r|n  (j�^  ]r}n  (h	he]r~n  (hh�e]rn  (hhe]r�n  (j�i  ]r�n  (h	h�e]r�n  (hh�eeee]r�n  (hhee]r�n  (h!]r�n  (h#h$e]r�n  (h	he]r�n  (hh�e]r�n  (h)heee]r�n  (j�^  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (h	h�e]r�n  (hh�e]r�n  (hhe]r�n  (j�^  ]r�n  (h	he]r�n  (hh�e]r�n  (hhe]r�n  (j�i  ]r�n  (h	h�e]r�n  (hh�eeee]r�n  (hhee]r�n  (h!]r�n  (h#h$e]r�n  (h	he]r�n  (hh�e]r�n  (h)heeej�n  j�n  j�n  j�n  j�n  j�n  j�n  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (h	h�e]r�n  (hh�e]r�n  (hhe]r�n  (j�^  ]r�n  (h	he]r�n  (hh�e]r�n  (hhe]r�n  (j�i  ]r�n  (h	h�e]r�n  (hh�eeee]r�n  (hhee]r�n  (h!]r�n  (h#h$e]r�n  (h	he]r�n  (hh�e]r�n  (h)heeej�n  j�n  j�n  j�n  j�n  j�n  j�n  j�n  j�n  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (h	h�e]r�n  (hh�e]r�n  (hhe]r�n  (j�^  ]r�n  (h	he]r�n  (hh�e]r�n  (hhe]r�n  (j�i  ]r�n  (h	h�e]r�n  (hh�eeee]r�n  (hhee]r�n  (h!]r�n  (h#h$e]r�n  (h	he]r�n  (hh�e]r�n  (h)heeej�n  j�n  j�n  j�n  j�n  j�n  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (h	h�e]r�n  (hh�e]r�n  (hhe]r�n  (j�^  ]r�n  (h	he]r�n  (hh�e]r�n  (hhe]r�n  (j�i  ]r�n  (h	h�e]r�n  (hh�eeee]r�n  (hhee]r�n  (h!]r�n  (h#h$e]r�n  (h	he]r�n  (hh�e]r�n  (h)heeej�n  j�n  j�n  j�n  j�n  j�n  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (h	h�e]r�n  (hh�e]r�n  (hhe]r�n  (j�^  ]r�n  (h	he]r�n  (hh�e]r�n  (hhe]r�n  (j�i  ]r�n  (h	h�e]r�n  (hh�eeee]r�n  (hhee]r�n  (h!]r�n  (h#h$e]r�n  (h	he]r�n  (hh�e]r�n  (h)heeej�n  j�n  j�n  j�n  j�n  j�n  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (h	h�e]r�n  (hh�e]r�n  (hhe]r�n  (j�^  ]r�n  (h	he]r�n  (hh�e]r�n  (hhe]r�n  (j�i  ]r�n  (h	h�e]r�n  (hh�eeee]r�n  (hhee]r�n  (h!]r�n  (h#h$e]r�n  (h	he]r�n  (hh�e]r�n  (h)heeej�n  j�n  j�n  j�n  j�n  j�n  j�n  j�n  j�n  j�n  j�n  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (j�^  ]r�n  (h	h�e]r�n  (hh�e]r o  (hhe]ro  (j�^  ]ro  (h	he]ro  (hh�e]ro  (hhe]ro  (j�i  ]ro  (h	h�e]ro  (hh�eeee]ro  (hhee]r	o  (h!]r
o  (h#h$e]ro  (h	he]ro  (hh�e]ro  (h)heeej�n  j�n  j�n  j�n  ]ro  (j�^  ]ro  (j�^  ]ro  (j�^  ]ro  (h	h�e]ro  (hh�e]ro  (hhe]ro  (j�^  ]ro  (h	he]ro  (hh�e]ro  (hhe]ro  (j�i  ]ro  (h	h�e]ro  (hh�eeee]ro  (hhee]ro  (h!]ro  (h#h$e]ro  (h	he]ro  (hh�e]r o  (h)heeejo  jo  jo  jo  jo  jo  jo  jo  jo  ]r!o  (j�^  ]r"o  (j�^  ]r#o  (j�^  ]r$o  (h	h�e]r%o  (hh�e]r&o  (hhe]r'o  (j�^  ]r(o  (h	he]r)o  (hh�e]r*o  (hhe]r+o  (j�i  ]r,o  (h	h�e]r-o  (hh�eeee]r.o  (hhee]r/o  (h!]r0o  (h#h$e]r1o  (h	he]r2o  (hh�e]r3o  (h)heeej!o  j!o  ]r4o  (j�^  ]r5o  (j�^  ]r6o  (j�^  ]r7o  (h	h�e]r8o  (hh�e]r9o  (hhe]r:o  (j�^  ]r;o  (h	he]r<o  (hh�e]r=o  (hhe]r>o  (j�i  ]r?o  (h	h�e]r@o  (hh�eeee]rAo  (hhee]rBo  (h!]rCo  (h#h$e]rDo  (h	he]rEo  (hh�e]rFo  (h)heeej4o  j4o  j4o  j4o  ]rGo  (j�^  ]rHo  (j�^  ]rIo  (j�^  ]rJo  (h	h�e]rKo  (hh�e]rLo  (hhe]rMo  (j�^  ]rNo  (h	he]rOo  (hh�e]rPo  (hhe]rQo  (j�i  ]rRo  (h	h�e]rSo  (hh�eeee]rTo  (hhee]rUo  (h!]rVo  (h#h$e]rWo  (h	he]rXo  (hh�e]rYo  (h)heee]rZo  (j�^  ]r[o  (j�^  ]r\o  (j�^  ]r]o  (h	h�e]r^o  (hh�e]r_o  (hhe]r`o  (j�^  ]rao  (h	he]rbo  (hh�e]rco  (hhe]rdo  (j�i  ]reo  (h	h�e]rfo  (hh�eeee]rgo  (hhee]rho  (h!]rio  (h#h$e]rjo  (h	he]rko  (hh�e]rlo  (h)heeejZo  jZo  ]rmo  (j�^  ]rno  (j�^  ]roo  (j�^  ]rpo  (h	h�e]rqo  (hh�e]rro  (hhe]rso  (j�^  ]rto  (h	he]ruo  (hh�e]rvo  (hhe]rwo  (j�i  ]rxo  (h	h�e]ryo  (hh�eeee]rzo  (hhee]r{o  (h!]r|o  (h#h$e]r}o  (h	he]r~o  (hh�e]ro  (h)heeejmo  jmo  jmo  jmo  ]r�o  (j�^  ]r�o  (j�^  ]r�o  (j�^  ]r�o  (h	h�e]r�o  (hh�e]r�o  (hhe]r�o  (j�^  ]r�o  (h	he]r�o  (hh�e]r�o  (hhe]r�o  (j�i  ]r�o  (h	h�e]r�o  (hh�eeee]r�o  (hhee]r�o  (h!]r�o  (h#h$e]r�o  (h	he]r�o  (hh�e]r�o  (h)heee]r�o  (j�^  ]r�o  (j�^  ]r�o  (j�^  ]r�o  (h	h�e]r�o  (hh�e]r�o  (hhe]r�o  (j�^  ]r�o  (h	he]r�o  (hh�e]r�o  (hhe]r�o  (j�i  ]r�o  (h	h�e]r�o  (hh�eeee]r�o  (hhee]r�o  (h!]r�o  (h#h$e]r�o  (h	he]r�o  (hh�e]r�o  (h)heeej�o  ]r�o  (j�^  ]r�o  (j�^  ]r�o  (j�^  ]r�o  (h	h�e]r�o  (hh�e]r�o  (hhe]r�o  (j�^  ]r�o  (h	he]r�o  (hh�e]r�o  (hhe]r�o  (j�i  ]r�o  (h	h�e]r�o  (hh�eeee]r�o  (hhee]r�o  (h!]r�o  (h#h$e]r�o  (h	he]r�o  (hh�e]r�o  (h)heee]r�o  (j�^  ]r�o  (j�^  ]r�o  (j�^  ]r�o  (h	h�e]r�o  (hh�e]r�o  (hhe]r�o  (j�^  ]r�o  (h	he]r�o  (hh�e]r�o  (hhe]r�o  (j�i  ]r�o  (h	h�e]r�o  (hh�eeee]r�o  (hhee]r�o  (h!]r�o  (h#h$e]r�o  (h	he]r�o  (hh�e]r�o  (h)heeej�o  j�o  ]r�o  (j�^  ]r�o  (j�^  ]r�o  (j�^  ]r�o  (h	h�e]r�o  (hh�e]r�o  (hhe]r�o  (j�^  ]r�o  (h	he]r�o  (hh�e]r�o  (hhe]r�o  (j�i  ]r�o  (h	h�e]r�o  (hh�eeee]r�o  (hhee]r�o  (h!]r�o  (h#h$e]r�o  (h	he]r�o  (hh�e]r�o  (h)heeej�o  j�o  ]r�o  (j�^  ]r�o  (j�^  ]r�o  (j�^  ]r�o  (h	h�e]r�o  (hh�e]r�o  (hhe]r�o  (j�^  ]r�o  (h	he]r�o  (hh�e]r�o  (hhe]r�o  (j�i  ]r�o  (h	h�e]r�o  (hh�eeee]r�o  (hhee]r�o  (h!]r�o  (h#h$e]r�o  (h	he]r�o  (hh�e]r�o  (h)heee]r�o  (j�^  ]r�o  (j�^  ]r�o  (j�^  ]r�o  (h	h�e]r�o  (hh�e]r�o  (hhe]r�o  (j�^  ]r�o  (h	he]r�o  (hh�e]r�o  (hhe]r�o  (j�i  ]r�o  (h	h�e]r�o  (hh�eeee]r�o  (hhee]r p  (h!]rp  (h#h$e]rp  (h	he]rp  (hh�e]rp  (h)heeej�o  j�o  j�o  j�o  ]rp  (j�^  ]rp  (j�^  ]rp  (j�^  ]rp  (h	h�e]r	p  (hh�e]r
p  (hhe]rp  (j�^  ]rp  (h	he]rp  (hh�e]rp  (hhe]rp  (j�i  ]rp  (h	h�e]rp  (hh�eeee]rp  (hhee]rp  (h!]rp  (h#h$e]rp  (h	he]rp  (hh�e]rp  (h)heee]rp  (j�^  ]rp  (j�^  ]rp  (j�^  ]rp  (h	h�e]rp  (hh�e]rp  (hhe]rp  (j�^  ]rp  (h	he]r p  (hh�e]r!p  (hhe]r"p  (j�i  ]r#p  (h	h�e]r$p  (hh�eeee]r%p  (hhee]r&p  (h!]r'p  (h#h$e]r(p  (h	he]r)p  (hh�e]r*p  (h)heeejp  jp  jp  ]r+p  (j�^  ]r,p  (j�^  ]r-p  (j�^  ]r.p  (h	h�e]r/p  (hh�e]r0p  (hhe]r1p  (j�^  ]r2p  (h	h�e]r3p  (hh�e]r4p  (hhe]r5p  (j�i  ]r6p  (h	h�e]r7p  (hh�eeee]r8p  (hhee]r9p  (h!]r:p  (h#h$e]r;p  (h	he]r<p  (hh�e]r=p  (h)heeej+p  j+p  ]r>p  (j�^  ]r?p  (j�^  ]r@p  (j�^  ]rAp  (h	h�e]rBp  (hh�e]rCp  (hhe]rDp  (j�^  ]rEp  (h	h�e]rFp  (hh�e]rGp  (hhe]rHp  (j�i  ]rIp  (h	h�e]rJp  (hh�eeee]rKp  (hhee]rLp  (h!]rMp  (h#h$e]rNp  (h	he]rOp  (hh�e]rPp  (h)heeej>p  j>p  ]rQp  (j�^  ]rRp  (j�^  ]rSp  (j�^  ]rTp  (h	h�e]rUp  (hh�e]rVp  (hhe]rWp  (j�^  ]rXp  (h	h�e]rYp  (hh�e]rZp  (hhe]r[p  (j�i  ]r\p  (h	h�e]r]p  (hh�eeee]r^p  (hhee]r_p  (h!]r`p  (h#h$e]rap  (h	he]rbp  (hh�e]rcp  (h)heeejQp  jQp  jQp  jQp  jQp  jQp  jQp  jQp  jQp  jQp  jQp  jQp  jQp  jQp  ]rdp  (j�^  ]rep  (j�^  ]rfp  (j�^  ]rgp  (h	h�e]rhp  (hh�e]rip  (hhe]rjp  (j�^  ]rkp  (h	h�e]rlp  (hh�e]rmp  (hhe]rnp  (j�i  ]rop  (h	h�e]rpp  (hh�eeee]rqp  (hhee]rrp  (h!]rsp  (h#h$e]rtp  (h	he]rup  (hh�e]rvp  (h)heeejdp  jdp  jdp  jdp  jdp  jdp  ]rwp  (j�^  ]rxp  (j�^  ]ryp  (j�^  ]rzp  (h	h�e]r{p  (hh�e]r|p  (hhe]r}p  (j�^  ]r~p  (h	h�e]rp  (hh�e]r�p  (hhe]r�p  (j�i  ]r�p  (h	h�e]r�p  (hh�eeee]r�p  (hhee]r�p  (h!]r�p  (h#h$e]r�p  (h	he]r�p  (hh�e]r�p  (h)heeejwp  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�i  ]r�p  (h	h�e]r�p  (hh�eeee]r�p  (hhee]r�p  (h!]r�p  (h#h$e]r�p  (h	he]r�p  (hh�e]r�p  (h)heee]r�p  (j�^  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�i  ]r�p  (h	h�e]r�p  (hh�eeee]r�p  (hhee]r�p  (h!]r�p  (h#h$e]r�p  (h	he]r�p  (hh�e]r�p  (h)heee]r�p  (j�^  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�i  ]r�p  (h	h�e]r�p  (hh�eeee]r�p  (hhee]r�p  (h!]r�p  (h#h$e]r�p  (h	he]r�p  (hh�e]r�p  (h)heeej�p  j�p  j�p  j�p  j�p  j�p  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�i  ]r�p  (h	h�e]r�p  (hh�eeee]r�p  (hhee]r�p  (h!]r�p  (h#h$e]r�p  (h	he]r�p  (hh�e]r�p  (h)heeej�p  j�p  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�i  ]r�p  (h	h�e]r�p  (hh�eeee]r�p  (hhee]r�p  (h!]r�p  (h#h$e]r�p  (h	he]r�p  (hh�e]r�p  (h)heeej�p  j�p  j�p  j�p  j�p  j�p  j�p  j�p  j�p  j�p  j�p  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�^  ]r�p  (h	h�e]r�p  (hh�e]r�p  (hhe]r�p  (j�i  ]r�p  (h	h�e]r�p  (hh�eeee]r�p  (hhee]r�p  (h!]r�p  (h#h$e]r�p  (h	he]r�p  (hh�e]r�p  (h)heeej�p  j�p  j�p  j�p  j�p  j�p  j�p  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (j�^  ]r�p  (h	h�e]r q  (hh�e]rq  (hhe]rq  (j�^  ]rq  (h	he]rq  (hh�e]rq  (hhe]rq  (j�i  ]rq  (h	h�e]rq  (hh�eeee]r	q  (hhee]r
q  (h!]rq  (h#h$e]rq  (h	he]rq  (hh�e]rq  (h)heee]rq  (j�^  ]rq  (j�^  ]rq  (j�^  ]rq  (h	h�e]rq  (hh�e]rq  (hhe]rq  (j�^  ]rq  (h	h�e]rq  (hh�e]rq  (hhe]rq  (j�i  ]rq  (h	h�e]rq  (hh�eeee]rq  (hhee]rq  (h!]rq  (h#h$e]rq  (h	he]r q  (hh�e]r!q  (h)heeejq  ]r"q  (j�^  ]r#q  (j�^  ]r$q  (j�^  ]r%q  (h	h�e]r&q  (hh�e]r'q  (hhe]r(q  (j�^  ]r)q  (h	h�e]r*q  (hh�e]r+q  (hhe]r,q  (j�i  ]r-q  (h	h�e]r.q  (hh�eeee]r/q  (hhee]r0q  (h!]r1q  (h#h$e]r2q  (h	he]r3q  (hh�e]r4q  (h)heeej"q  j"q  j"q  j"q  j"q  j"q  ]r5q  (j�^  ]r6q  (j�^  ]r7q  (j�^  ]r8q  (h	h�e]r9q  (hh�e]r:q  (hhe]r;q  (j�^  ]r<q  (h	h�e]r=q  (hh�e]r>q  (hhe]r?q  (j�i  ]r@q  (h	h�e]rAq  (hh�eeee]rBq  (hhee]rCq  (h!]rDq  (h#h$e]rEq  (h	he]rFq  (hh�e]rGq  (h)heeej5q  j5q  j5q  j5q  j5q  ]rHq  (j�^  ]rIq  (j�^  ]rJq  (j�^  ]rKq  (h	h�e]rLq  (hh�e]rMq  (hhe]rNq  (j�^  ]rOq  (h	h�e]rPq  (hh�e]rQq  (hhe]rRq  (j�i  ]rSq  (h	h�e]rTq  (hh�eeee]rUq  (hhee]rVq  (h!]rWq  (h#h$e]rXq  (h	he]rYq  (hh�e]rZq  (h)heeejHq  jHq  ]r[q  (j�^  ]r\q  (j�^  ]r]q  (j�^  ]r^q  (h	h�e]r_q  (hh�e]r`q  (hhe]raq  (j�^  ]rbq  (h	h�e]rcq  (hh�e]rdq  (hhe]req  (j�i  ]rfq  (h	h�e]rgq  (hh�eeee]rhq  (hhee]riq  (h!]rjq  (h#h$e]rkq  (h	he]rlq  (hh�e]rmq  (h)heee]rnq  (j�^  ]roq  (j�^  ]rpq  (j�^  ]rqq  (h	h�e]rrq  (hh�e]rsq  (hhe]rtq  (j�^  ]ruq  (h	h�e]rvq  (hh�e]rwq  (hhe]rxq  (j�i  ]ryq  (h	h�e]rzq  (hh�eeee]r{q  (hhee]r|q  (h!]r}q  (h#h$e]r~q  (h	he]rq  (hh�e]r�q  (h)heee]r�q  (j�^  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�i  ]r�q  (h	h�e]r�q  (hh�eeee]r�q  (hhee]r�q  (h!]r�q  (h#h$e]r�q  (h	he]r�q  (hh�e]r�q  (h)heeej�q  j�q  j�q  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�i  ]r�q  (h	h�e]r�q  (hh�eeee]r�q  (hhee]r�q  (h!]r�q  (h#h$e]r�q  (h	he]r�q  (hh�e]r�q  (h)heeej�q  j�q  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�i  ]r�q  (h	h�e]r�q  (hh�eeee]r�q  (hhee]r�q  (h!]r�q  (h#h$e]r�q  (h	he]r�q  (hh�e]r�q  (h)heeej�q  j�q  j�q  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�i  ]r�q  (h	h�e]r�q  (hh�eeee]r�q  (hhee]r�q  (h!]r�q  (h#h$e]r�q  (h	he]r�q  (hh�e]r�q  (h)heee]r�q  (j�^  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�i  ]r�q  (h	h�e]r�q  (hh�eeee]r�q  (hhee]r�q  (h!]r�q  (h#h$e]r�q  (h	he]r�q  (hh�e]r�q  (h)heeej�q  j�q  j�q  j�q  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�^  ]r�q  (h	he]r�q  (hh�e]r�q  (hhe]r�q  (j�i  ]r�q  (h	h�e]r�q  (hh�eeee]r�q  (hhee]r�q  (h!]r�q  (h#h$e]r�q  (h	he]r�q  (hh�e]r�q  (h)heeej�q  j�q  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (j�^  ]r�q  (h	h�e]r�q  (hh�e]r�q  (hhe]r�q  (j�^  ]r�q  (h	he]r�q  (hh�e]r�q  (hhe]r�q  (j�i  ]r�q  (h	h�e]r�q  (hh�eeee]r r  (hhee]rr  (h!]rr  (h#h$e]rr  (h	he]rr  (hh�e]rr  (h)heeej�q  j�q  j�q  ]rr  (j�^  ]rr  (j�^  ]rr  (j�^  ]r	r  (h	h�e]r
r  (hh�e]rr  (hhe]rr  (j�^  ]rr  (h	he]rr  (hh�e]rr  (hhe]rr  (j�i  ]rr  (h	h�e]rr  (hh�eeee]rr  (hhee]rr  (h!]rr  (h#h$e]rr  (h	he]rr  (hh�e]rr  (h)heeejr  ]rr  (j�^  ]rr  (j�^  ]rr  (j�^  ]rr  (h	h�e]rr  (hh�e]rr  (hhe]rr  (j�^  ]r r  (h	he]r!r  (hh�e]r"r  (hhe]r#r  (j�i  ]r$r  (h	h�e]r%r  (hh�eeee]r&r  (hhee]r'r  (h!]r(r  (h#h$e]r)r  (h	he]r*r  (hh�e]r+r  (h)heee]r,r  (j�^  ]r-r  (j�^  ]r.r  (j�^  ]r/r  (h	h�e]r0r  (hh�e]r1r  (hhe]r2r  (j�^  ]r3r  (h	he]r4r  (hh�e]r5r  (hhe]r6r  (j�i  ]r7r  (h	h�e]r8r  (hh�eeee]r9r  (hhee]r:r  (h!]r;r  (h#h$e]r<r  (h	he]r=r  (hh�e]r>r  (h)heee]r?r  (j�^  ]r@r  (j�^  ]rAr  (j�^  ]rBr  (h	h�e]rCr  (hh�e]rDr  (hhe]rEr  (j�^  ]rFr  (h	he]rGr  (hh�e]rHr  (hhe]rIr  (j�i  ]rJr  (h	h�e]rKr  (hh�eeee]rLr  (hhee]rMr  (h!]rNr  (h#h$e]rOr  (h	he]rPr  (hh�e]rQr  (h)heeej?r  j?r  j?r  j?r  ]rRr  (j�^  ]rSr  (j�^  ]rTr  (j�^  ]rUr  (h	h�e]rVr  (hh�e]rWr  (hhe]rXr  (j�^  ]rYr  (h	he]rZr  (hh�e]r[r  (hhe]r\r  (j�i  ]r]r  (h	h�e]r^r  (hh�eeee]r_r  (hhee]r`r  (h!]rar  (h#h$e]rbr  (h	he]rcr  (hh�e]rdr  (h)heeejRr  jRr  jRr  jRr  ]rer  (j�^  ]rfr  (j�^  ]rgr  (j�^  ]rhr  (h	h�e]rir  (hh�e]rjr  (hhe]rkr  (j�^  ]rlr  (h	he]rmr  (hh�e]rnr  (hhe]ror  (j�i  ]rpr  (h	h�e]rqr  (hh�eeee]rrr  (hhee]rsr  (h!]rtr  (h#h$e]rur  (h	he]rvr  (hh�e]rwr  (h)heeejer  jer  ]rxr  (j�^  ]ryr  (j�^  ]rzr  (j�^  ]r{r  (h	h�e]r|r  (hh�e]r}r  (hhe]r~r  (j�^  ]rr  (h	he]r�r  (hh�e]r�r  (hhe]r�r  (j�i  ]r�r  (h	h�e]r�r  (hh�eeee]r�r  (hhee]r�r  (h!]r�r  (h#h$e]r�r  (h	he]r�r  (hh�e]r�r  (h)heeejxr  ]r�r  (j�^  ]r�r  (j�^  ]r�r  (j�^  ]r�r  (h	h�e]r�r  (hh�e]r�r  (hhe]r�r  (j�^  ]r�r  (h	he]r�r  (hh�e]r�r  (hhe]r�r  (j�i  ]r�r  (h	h�e]r�r  (hh�eeee]r�r  (hhee]r�r  (h!]r�r  (h#h$e]r�r  (h	he]r�r  (hh�e]r�r  (h)heeej�r  j�r  ]r�r  (j�^  ]r�r  (j�^  ]r�r  (j�^  ]r�r  (h	h�e]r�r  (hh�e]r�r  (hhe]r�r  (j�^  ]r�r  (h	he]r�r  (hh�e]r�r  (hhe]r�r  (j�i  ]r�r  (h	h�e]r�r  (hh�eeee]r�r  (hhee]r�r  (h!]r�r  (h#h$e]r�r  (h	he]r�r  (hh�e]r�r  (h)heeej�r  j�r  j�r  j�r  j�r  j�r  j�r  j�r  ]r�r  (j�^  ]r�r  (j�^  ]r�r  (j�^  ]r�r  (h	h�e]r�r  (hh�e]r�r  (hhe]r�r  (j�^  ]r�r  (h	h�e]r�r  (hh�e]r�r  (hhe]r�r  (j�i  ]r�r  (h	h�e]r�r  (hh�eeee]r�r  (hhee]r�r  (h!]r�r  (h#h$e]r�r  (h	he]r�r  (hh�e]r�r  (h)heee]r�r  (j�^  ]r�r  (j�^  ]r�r  (j�^  ]r�r  (h	h�e]r�r  (hh�e]r�r  (hhe]r�r  (j�^  ]r�r  (h	h�e]r�r  (hh�e]r�r  (hhe]r�r  (j�i  ]r�r  (h	h�e]r�r  (hh�eeee]r�r  (hhee]r�r  (h!]r�r  (h#h$e]r�r  (h	he]r�r  (hh�e]r�r  (h)heeej�r  ]r�r  (j�^  ]r�r  (j�^  ]r�r  (j�^  ]r�r  (h	h�e]r�r  (hh�e]r�r  (hhe]r�r  (j�^  ]r�r  (h	he]r�r  (hh�e]r�r  (hhe]r�r  (j�i  ]r�r  (h	h�e]r�r  (hh�eeee]r�r  (hhee]r�r  (h!]r�r  (h#h$e]r�r  (h	he]r�r  (hh�e]r�r  (h)heeej�r  j�r  j�r  j�r  j�r  ]r�r  (j�^  ]r�r  (j�^  ]r�r  (j�^  ]r�r  (h	h�e]r�r  (hh�e]r�r  (hhe]r�r  (j�^  ]r�r  (h	he]r�r  (hh�e]r�r  (hhe]r�r  (j�i  ]r�r  (h	h�e]r�r  (hh�eeee]r�r  (hhee]r�r  (h!]r�r  (h#h$e]r�r  (h	he]r�r  (hh�e]r�r  (h)heee]r�r  (j�^  ]r�r  (j�^  ]r�r  (j�^  ]r s  (h	h�e]rs  (hh�e]rs  (hhe]rs  (j�^  ]rs  (h	he]rs  (hh�e]rs  (hhe]rs  (j�i  ]rs  (h	h�e]r	s  (hh�eeee]r
s  (hhee]rs  (h!]rs  (h#h$e]rs  (h	he]rs  (hh�e]rs  (h)heeej�r  ]rs  (j�^  ]rs  (j�^  ]rs  (j�^  ]rs  (h	h�e]rs  (hh�e]rs  (hhe]rs  (j�^  ]rs  (h	he]rs  (hh�e]rs  (hhe]rs  (j�i  ]rs  (h	h�e]rs  (hh�eeee]rs  (hhee]rs  (h!]rs  (h#h$e]r s  (h	he]r!s  (hh�e]r"s  (h)heeejs  js  js  ]r#s  (j�^  ]r$s  (j�^  ]r%s  (j�^  ]r&s  (h	h�e]r's  (hh�e]r(s  (hhe]r)s  (j�^  ]r*s  (h	h�e]r+s  (hh�e]r,s  (hhe]r-s  (j�i  ]r.s  (h	h�e]r/s  (hh�eeee]r0s  (hhee]r1s  (h!]r2s  (h#h$e]r3s  (h	he]r4s  (hh�e]r5s  (h)heeej#s  j#s  j#s  j#s  ]r6s  (j�^  ]r7s  (j�^  ]r8s  (j�^  ]r9s  (h	h�e]r:s  (hh�e]r;s  (hhe]r<s  (j�^  ]r=s  (h	h�e]r>s  (hh�e]r?s  (hhe]r@s  (j�i  ]rAs  (h	h�e]rBs  (hh�eeee]rCs  (hhee]rDs  (h!]rEs  (h#h$e]rFs  (h	he]rGs  (hh�e]rHs  (h)heeej6s  ]rIs  (j�^  ]rJs  (j�^  ]rKs  (j�^  ]rLs  (h	h�e]rMs  (hh�e]rNs  (hhe]rOs  (j�^  ]rPs  (h	h�e]rQs  (hh�e]rRs  (hhe]rSs  (j�i  ]rTs  (h	h�e]rUs  (hh�eeee]rVs  (hhee]rWs  (h!]rXs  (h#h$e]rYs  (h	he]rZs  (hh�e]r[s  (h)heeejIs  ]r\s  (j�^  ]r]s  (j�^  ]r^s  (j�^  ]r_s  (h	h�e]r`s  (hh�e]ras  (hhe]rbs  (j�^  ]rcs  (h	he]rds  (hh�e]res  (hhe]rfs  (j�i  ]rgs  (h	h�e]rhs  (hh�eeee]ris  (hhee]rjs  (h!]rks  (h#h$e]rls  (h	he]rms  (hh�e]rns  (h)heeej\s  j\s  j\s  j\s  j\s  ]ros  (j�^  ]rps  (j�^  ]rqs  (j�^  ]rrs  (h	h�e]rss  (hh�e]rts  (hhe]rus  (j�^  ]rvs  (h	he]rws  (hh�e]rxs  (hhe]rys  (j�i  ]rzs  (h	h�e]r{s  (hh�eeee]r|s  (hhee]r}s  (h!]r~s  (h#h$e]rs  (h	he]r�s  (hh�e]r�s  (h)heee]r�s  (j�^  ]r�s  (j�^  ]r�s  (j�^  ]r�s  (h	h�e]r�s  (hh�e]r�s  (hhe]r�s  (j�^  ]r�s  (h	he]r�s  (hh�e]r�s  (hhe]r�s  (X	   Next-Mover�s  ]r�s  (h	h�e]r�s  (hh�eeee]r�s  (hhee]r�s  (h!]r�s  (h#h$e]r�s  (h	he]r�s  (hh�e]r�s  (h)heee]r�s  (j�^  ]r�s  (j�^  ]r�s  (j�^  ]r�s  (h	h�e]r�s  (hh�e]r�s  (hhe]r�s  (j�^  ]r�s  (h	he]r�s  (hh�e]r�s  (hhe]r�s  (j�s  ]r�s  (h	h�e]r�s  (hh�eeee]r�s  (hhee]r�s  (h!]r�s  (h#h$e]r�s  (h	he]r�s  (hh�e]r�s  (h)heeej�s  ]r�s  (j�^  ]r�s  (j�^  ]r�s  (j�^  ]r�s  (h	h�e]r�s  (hh�e]r�s  (hhe]r�s  (j�^  ]r�s  (h	he]r�s  (hh�e]r�s  (hhe]r�s  (j�s  ]r�s  (h	h�e]r�s  (hh�eeee]r�s  (hhee]r�s  (h!]r�s  (h#h$e]r�s  (h	he]r�s  (hh�e]r�s  (h)heee]r�s  (j�^  ]r�s  (j�^  ]r�s  (j�^  ]r�s  (h	h�e]r�s  (hh�e]r�s  (hhe]r�s  (j�^  ]r�s  (h	he]r�s  (hh�e]r�s  (hhe]r�s  (j�s  ]r�s  (h	h�e]r�s  (hh�eeee]r�s  (hhee]r�s  (h!]r�s  (h#h$e]r�s  (h	he]r�s  (hh�e]r�s  (h)heeej�s  j�s  j�s  j�s  j�s  ]r�s  (j�^  ]r�s  (j�^  ]r�s  (j�^  ]r�s  (h	h�e]r�s  (hh�e]r�s  (hhe]r�s  (j�^  ]r�s  (h	he]r�s  (hh�e]r�s  (hhe]r�s  (j�s  ]r�s  (h	h�e]r�s  (hh�eeee]r�s  (hhee]r�s  (h!]r�s  (h#h$e]r�s  (h	he]r�s  (hh�e]r�s  (h)heeej�s  j�s  ]r�s  (j�^  ]r�s  (j�^  ]r�s  (j�^  ]r�s  (h	h�e]r�s  (hh�e]r�s  (hhe]r�s  (j�^  ]r�s  (h	he]r�s  (hh�e]r�s  (hhe]r�s  (j�s  ]r�s  (h	h�e]r�s  (hh�eeee]r�s  (hhee]r�s  (h!]r�s  (h#h$e]r�s  (h	he]r�s  (hh�e]r�s  (h)heeej�s  ]r�s  (j�^  ]r�s  (j�^  ]r�s  (j�^  ]r�s  (h	h�e]r�s  (hh�e]r�s  (hhe]r�s  (j�^  ]r�s  (h	he]r�s  (hh�e]r�s  (hhe]r�s  (j�s  ]r t  (h	h�e]rt  (hh�eeee]rt  (hhee]rt  (h!]rt  (h#h$e]rt  (h	he]rt  (hh�e]rt  (h)heeej�s  j�s  j�s  j�s  j�s  j�s  j�s  j�s  ]rt  (j�^  ]r	t  (j�^  ]r
t  (j�^  ]rt  (h	h�e]rt  (hh�e]rt  (hhe]rt  (j�^  ]rt  (h	he]rt  (hh�e]rt  (hhe]rt  (j�s  ]rt  (h	h�e]rt  (hh�eeee]rt  (hhee]rt  (h!]rt  (h#h$e]rt  (h	he]rt  (hh�e]rt  (h)heeejt  ]rt  (j�^  ]rt  (j�^  ]rt  (j�^  ]rt  (h	h�e]rt  (hh�e]r t  (hhe]r!t  (j�^  ]r"t  (h	he]r#t  (hh�e]r$t  (hhe]r%t  (j�s  ]r&t  (h	h�e]r't  (hh�eeee]r(t  (hhee]r)t  (h!]r*t  (h#h$e]r+t  (h	he]r,t  (hh�e]r-t  (h)heeejt  jt  jt  jt  jt  jt  jt  ]r.t  (j�^  ]r/t  (j�^  ]r0t  (j�^  ]r1t  (h	h�e]r2t  (hh�e]r3t  (hhe]r4t  (j�^  ]r5t  (h	he]r6t  (hh�e]r7t  (hhe]r8t  (j�s  ]r9t  (h	h�e]r:t  (hh�eeee]r;t  (hhee]r<t  (h!]r=t  (h#h$e]r>t  (h	he]r?t  (hh�e]r@t  (h)heeej.t  j.t  j.t  j.t  j.t  j.t  j.t  ]rAt  (j�^  ]rBt  (j�^  ]rCt  (j�^  ]rDt  (h	h�e]rEt  (hh�e]rFt  (hhe]rGt  (j�^  ]rHt  (h	h�e]rIt  (hh�e]rJt  (hhe]rKt  (j�s  ]rLt  (h	h�e]rMt  (hh�eeee]rNt  (hhee]rOt  (h!]rPt  (h#h$e]rQt  (h	he]rRt  (hh�e]rSt  (h)heeejAt  jAt  jAt  ]rTt  (j�^  ]rUt  (j�^  ]rVt  (j�^  ]rWt  (h	h�e]rXt  (hh�e]rYt  (hhe]rZt  (j�^  ]r[t  (h	h�e]r\t  (hh�e]r]t  (hhe]r^t  (j�s  ]r_t  (h	h�e]r`t  (hh�eeee]rat  (hhee]rbt  (h!]rct  (h#h$e]rdt  (h	he]ret  (hh�e]rft  (h)heeejTt  jTt  jTt  jTt  jTt  jTt  jTt  jTt  jTt  jTt  jTt  jTt  jTt  jTt  jTt  jTt  ]rgt  (j�^  ]rht  (j�^  ]rit  (j�^  ]rjt  (h	h�e]rkt  (hh�e]rlt  (hhe]rmt  (j�^  ]rnt  (h	h�e]rot  (hh�e]rpt  (hhe]rqt  (j�s  ]rrt  (h	h�e]rst  (hh�eeee]rtt  (hhee]rut  (h!]rvt  (h#h$e]rwt  (h	he]rxt  (hh�e]ryt  (h)heeejgt  e(jgt  jgt  jgt  jgt  jgt  jgt  jgt  jgt  jgt  jgt  ]rzt  (j�^  ]r{t  (j�^  ]r|t  (j�^  ]r}t  (h	h�e]r~t  (hh�e]rt  (hhe]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�s  ]r�t  (h	h�e]r�t  (hh�eeee]r�t  (hhee]r�t  (h!]r�t  (h#h$e]r�t  (h	he]r�t  (hh�e]r�t  (h)heee]r�t  (j�^  ]r�t  (j�^  ]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�s  ]r�t  (h	h�e]r�t  (hh�eeee]r�t  (hhee]r�t  (h!]r�t  (h#h$e]r�t  (h	he]r�t  (hh�e]r�t  (h)heeej�t  j�t  j�t  j�t  ]r�t  (j�^  ]r�t  (j�^  ]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�s  ]r�t  (h	h�e]r�t  (hh�eeee]r�t  (hhee]r�t  (h!]r�t  (h#h$e]r�t  (h	he]r�t  (hh�e]r�t  (h)heeej�t  j�t  j�t  j�t  j�t  j�t  j�t  ]r�t  (j�^  ]r�t  (j�^  ]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�s  ]r�t  (h	h�e]r�t  (hh�eeee]r�t  (hhee]r�t  (h!]r�t  (h#h$e]r�t  (h	he]r�t  (hh�e]r�t  (h)heee]r�t  (j�^  ]r�t  (j�^  ]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�s  ]r�t  (h	h�e]r�t  (hh�eeee]r�t  (hhee]r�t  (h!]r�t  (h#h$e]r�t  (h	he]r�t  (hh�e]r�t  (h)heeej�t  j�t  ]r�t  (j�^  ]r�t  (j�^  ]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�s  ]r�t  (h	h�e]r�t  (hh�eeee]r�t  (hhee]r�t  (h!]r�t  (h#h$e]r�t  (h	he]r�t  (hh�e]r�t  (h)heee]r�t  (j�^  ]r�t  (j�^  ]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�^  ]r�t  (h	h�e]r�t  (hh�e]r�t  (hhe]r�t  (j�s  ]r�t  (h	h�e]r�t  (hh�eeee]r�t  (hhee]r�t  (h!]r�t  (h#h$e]r�t  (h	he]r�t  (hh�e]r�t  (h)heee]r�t  (j�^  ]r u  (j�^  ]ru  (j�^  ]ru  (h	h�e]ru  (hh�e]ru  (hhe]ru  (j�^  ]ru  (h	h�e]ru  (hh�e]ru  (hhe]r	u  (j�s  ]r
u  (h	h�e]ru  (hh�eeee]ru  (hhee]ru  (h!]ru  (h#h$e]ru  (h	he]ru  (hh�e]ru  (h)heeej�t  j�t  ]ru  (j�^  ]ru  (j�^  ]ru  (j�^  ]ru  (h	h�e]ru  (hh�e]ru  (hhe]ru  (j�^  ]ru  (h	h�e]ru  (hh�e]ru  (hhe]ru  (j�s  ]ru  (h	h�e]ru  (hh�eeee]ru  (hhee]r u  (h!]r!u  (h#h$e]r"u  (h	he]r#u  (hh�e]r$u  (h)heeeju  ju  ju  ju  ju  ju  ju  ju  ju  ju  ju  ju  ]r%u  (j�^  ]r&u  (j�^  ]r'u  (j�^  ]r(u  (h	h�e]r)u  (hh�e]r*u  (hhe]r+u  (j�^  ]r,u  (h	h�e]r-u  (hh�e]r.u  (hhe]r/u  (j�s  ]r0u  (h	h�e]r1u  (hh�eeee]r2u  (hhee]r3u  (h!]r4u  (h#h$e]r5u  (h	he]r6u  (hh�e]r7u  (h)heeej%u  j%u  j%u  j%u  j%u  j%u  j%u  j%u  j%u  ]r8u  (j�^  ]r9u  (j�^  ]r:u  (j�^  ]r;u  (h	h�e]r<u  (hh�e]r=u  (hhe]r>u  (j�^  ]r?u  (h	h�e]r@u  (hh�e]rAu  (hhe]rBu  (j�s  ]rCu  (h	h�e]rDu  (hh�eeee]rEu  (hhee]rFu  (h!]rGu  (h#h$e]rHu  (h	he]rIu  (hh�e]rJu  (h)heeej8u  j8u  j8u  j8u  j8u  j8u  ]rKu  (j�^  ]rLu  (j�^  ]rMu  (j�^  ]rNu  (h	h�e]rOu  (hh�e]rPu  (hhe]rQu  (j�^  ]rRu  (h	h�e]rSu  (hh�e]rTu  (hhe]rUu  (j�s  ]rVu  (h	h�e]rWu  (hh�eeee]rXu  (hhee]rYu  (h!]rZu  (h#h$e]r[u  (h	he]r\u  (hh�e]r]u  (h)heeejKu  ]r^u  (j�^  ]r_u  (j�^  ]r`u  (j�^  ]rau  (h	h�e]rbu  (hh�e]rcu  (hhe]rdu  (j�^  ]reu  (h	he]rfu  (hh�e]rgu  (hhe]rhu  (j�s  ]riu  (h	h�e]rju  (hh�eeee]rku  (hhee]rlu  (h!]rmu  (h#h$e]rnu  (h	he]rou  (hh�e]rpu  (h)heeej^u  j^u  j^u  j^u  j^u  j^u  j^u  j^u  j^u  j^u  ]rqu  (j�^  ]rru  (j�^  ]rsu  (j�^  ]rtu  (h	h�e]ruu  (hh�e]rvu  (hhe]rwu  (j�^  ]rxu  (h	he]ryu  (hh�e]rzu  (hhe]r{u  (j�s  ]r|u  (h	h�e]r}u  (hh�eeee]r~u  (hhee]ru  (h!]r�u  (h#h$e]r�u  (h	he]r�u  (hh�e]r�u  (h)heeejqu  jqu  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (h	h�e]r�u  (hh�e]r�u  (hhe]r�u  (j�^  ]r�u  (h	he]r�u  (hh�e]r�u  (hhe]r�u  (j�s  ]r�u  (h	h�e]r�u  (hh�eeee]r�u  (hhee]r�u  (h!]r�u  (h#h$e]r�u  (h	he]r�u  (hh�e]r�u  (h)heee]r�u  (j�^  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (h	h�e]r�u  (hh�e]r�u  (hhe]r�u  (j�^  ]r�u  (h	he]r�u  (hh�e]r�u  (hhe]r�u  (j�s  ]r�u  (h	h�e]r�u  (hh�eeee]r�u  (hhee]r�u  (h!]r�u  (h#h$e]r�u  (h	he]r�u  (hh�e]r�u  (h)heeej�u  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (h	h�e]r�u  (hh�e]r�u  (hhe]r�u  (j�^  ]r�u  (h	he]r�u  (hh�e]r�u  (hhe]r�u  (j�s  ]r�u  (h	h�e]r�u  (hh�eeee]r�u  (hhee]r�u  (h!]r�u  (h#h$e]r�u  (h	he]r�u  (hh�e]r�u  (h)heeej�u  j�u  j�u  j�u  j�u  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (h	h�e]r�u  (hh�e]r�u  (hhe]r�u  (j�^  ]r�u  (h	he]r�u  (hh�e]r�u  (hhe]r�u  (j�s  ]r�u  (h	h�e]r�u  (hh�eeee]r�u  (hhee]r�u  (h!]r�u  (h#h$e]r�u  (h	he]r�u  (hh�e]r�u  (h)heeej�u  j�u  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (h	h�e]r�u  (hh�e]r�u  (hhe]r�u  (j�^  ]r�u  (h	he]r�u  (hh�e]r�u  (hhe]r�u  (j�s  ]r�u  (h	h�e]r�u  (hh�eeee]r�u  (hhee]r�u  (h!]r�u  (h#h$e]r�u  (h	he]r�u  (hh�e]r�u  (h)heeej�u  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (h	h�e]r�u  (hh�e]r�u  (hhe]r�u  (j�^  ]r�u  (h	he]r�u  (hh�e]r�u  (hhe]r�u  (j�s  ]r�u  (h	h�e]r�u  (hh�eeee]r�u  (hhee]r�u  (h!]r�u  (h#h$e]r�u  (h	he]r�u  (hh�e]r�u  (h)heee]r�u  (j�^  ]r�u  (j�^  ]r�u  (j�^  ]r�u  (h	h�e]r�u  (hh�e]r�u  (hhe]r�u  (j�^  ]r�u  (h	he]r�u  (hh�e]r�u  (hhe]r v  (j�s  ]rv  (h	h�e]rv  (hh�eeee]rv  (hhee]rv  (h!]rv  (h#h$e]rv  (h	he]rv  (hh�e]rv  (h)heeej�u  j�u  ]r	v  (j�^  ]r
v  (j�^  ]rv  (j�^  ]rv  (h	h�e]rv  (hh�e]rv  (hhe]rv  (j�^  ]rv  (h	he]rv  (hh�e]rv  (hhe]rv  (j�s  ]rv  (h	h�e]rv  (hh�eeee]rv  (hhee]rv  (h!]rv  (h#h$e]rv  (h	he]rv  (hh�e]rv  (h)heeej	v  j	v  j	v  j	v  j	v  j	v  j	v  j	v  j	v  j	v  j	v  j	v  j	v  j	v  j	v  j	v  j	v  ]rv  (j�^  ]rv  (j�^  ]rv  (j�^  ]rv  (h	h�e]r v  (hh�e]r!v  (hhe]r"v  (j�^  ]r#v  (h	he]r$v  (hh�e]r%v  (hhe]r&v  (j�s  ]r'v  (h	h�e]r(v  (hh�eeee]r)v  (hhee]r*v  (h!]r+v  (h#h$e]r,v  (h	he]r-v  (hh�e]r.v  (h)heee]r/v  (j�^  ]r0v  (j�^  ]r1v  (j�^  ]r2v  (h	h�e]r3v  (hh�e]r4v  (hhe]r5v  (j�^  ]r6v  (h	he]r7v  (hh�e]r8v  (hhe]r9v  (j�s  ]r:v  (h	h�e]r;v  (hh�eeee]r<v  (hhee]r=v  (h!]r>v  (h#h$e]r?v  (h	he]r@v  (hh�e]rAv  (h)heeej/v  ]rBv  (j�^  ]rCv  (j�^  ]rDv  (j�^  ]rEv  (h	h�e]rFv  (hh�e]rGv  (hhe]rHv  (j�^  ]rIv  (h	he]rJv  (hh�e]rKv  (hhe]rLv  (j�s  ]rMv  (h	h�e]rNv  (hh�eeee]rOv  (hhee]rPv  (h!]rQv  (h#h$e]rRv  (h	he]rSv  (hh�e]rTv  (h)heee]rUv  (j�^  ]rVv  (j�^  ]rWv  (j�^  ]rXv  (h	h�e]rYv  (hh�e]rZv  (hhe]r[v  (j�^  ]r\v  (h	he]r]v  (hh�e]r^v  (hhe]r_v  (j�s  ]r`v  (h	h�e]rav  (hh�eeee]rbv  (hhee]rcv  (h!]rdv  (h#h$e]rev  (h	he]rfv  (hh�e]rgv  (h)heeejUv  jUv  jUv  ]rhv  (j�^  ]riv  (j�^  ]rjv  (j�^  ]rkv  (h	h�e]rlv  (hh�e]rmv  (hhe]rnv  (j�^  ]rov  (h	he]rpv  (hh�e]rqv  (hhe]rrv  (j�s  ]rsv  (h	h�e]rtv  (hh�eeee]ruv  (hhee]rvv  (h!]rwv  (h#h$e]rxv  (h	he]ryv  (hh�e]rzv  (h)heeejhv  jhv  jhv  ]r{v  (j�^  ]r|v  (j�^  ]r}v  (j�^  ]r~v  (h	h�e]rv  (hh�e]r�v  (hhe]r�v  (j�^  ]r�v  (h	he]r�v  (hh�e]r�v  (hhe]r�v  (j�s  ]r�v  (h	h�e]r�v  (hh�eeee]r�v  (hhee]r�v  (h!]r�v  (h#h$e]r�v  (h	he]r�v  (hh�e]r�v  (h)heeej{v  ]r�v  (j�^  ]r�v  (j�^  ]r�v  (j�^  ]r�v  (h	h�e]r�v  (hh�e]r�v  (hhe]r�v  (j�^  ]r�v  (h	he]r�v  (hh�e]r�v  (hhe]r�v  (j�s  ]r�v  (h	h�e]r�v  (hh�eeee]r�v  (hhee]r�v  (h!]r�v  (h#h$e]r�v  (h	he]r�v  (hh�e]r�v  (h)heeej�v  ]r�v  (j�^  ]r�v  (j�^  ]r�v  (j�^  ]r�v  (h	h�e]r�v  (hh�e]r�v  (hhe]r�v  (j�^  ]r�v  (h	he]r�v  (hh�e]r�v  (hhe]r�v  (j�s  ]r�v  (h	h�e]r�v  (hh�eeee]r�v  (hhee]r�v  (h!]r�v  (h#h$e]r�v  (h	he]r�v  (hh�e]r�v  (h)heeej�v  j�v  j�v  ]r�v  (j�^  ]r�v  (j�^  ]r�v  (j�^  ]r�v  (h	h�e]r�v  (hh�e]r�v  (hhe]r�v  (j�^  ]r�v  (h	he]r�v  (hh�e]r�v  (hhe]r�v  (j�s  ]r�v  (h	h�e]r�v  (hh�eeee]r�v  (hhee]r�v  (h!]r�v  (h#h$e]r�v  (h	he]r�v  (hh�e]r�v  (h)heeej�v  j�v  ]r�v  (j�^  ]r�v  (j�^  ]r�v  (j�^  ]r�v  (h	h�e]r�v  (hh�e]r�v  (hhe]r�v  (j�^  ]r�v  (h	he]r�v  (hh�e]r�v  (hhe]r�v  (j�s  ]r�v  (h	h�e]r�v  (hh�eeee]r�v  (hhee]r�v  (h!]r�v  (h#h$e]r�v  (h	he]r�v  (hh�e]r�v  (h)heeej�v  j�v  j�v  j�v  j�v  j�v  j�v  j�v  j�v  ]r�v  (j�^  ]r�v  (j�^  ]r�v  (j�^  ]r�v  (h	h�e]r�v  (hh�e]r�v  (hhe]r�v  (j�^  ]r�v  (h	he]r�v  (hh�e]r�v  (hhe]r�v  (j�s  ]r�v  (h	h�e]r�v  (hh�eeee]r�v  (hhee]r�v  (h!]r�v  (h#h$e]r�v  (h	he]r�v  (hh�e]r�v  (h)heee]r�v  (j�^  ]r�v  (j�^  ]r�v  (j�^  ]r�v  (h	h�e]r�v  (hh�e]r�v  (hhe]r�v  (j�^  ]r�v  (h	he]r�v  (hh�e]r�v  (hhe]r�v  (j�s  ]r�v  (h	h�e]r�v  (hh�eeee]r�v  (hhee]r�v  (h!]r�v  (h#h$e]r�v  (h	he]r�v  (hh�e]r�v  (h)heee]r w  (j�^  ]rw  (j�^  ]rw  (j�^  ]rw  (h	h�e]rw  (hh�e]rw  (hhe]rw  (j�^  ]rw  (h	he]rw  (hh�e]r	w  (hhe]r
w  (j�s  ]rw  (h	h�e]rw  (hh�eeee]rw  (hhee]rw  (h!]rw  (h#h$e]rw  (h	he]rw  (hh�e]rw  (h)heeej w  j w  ]rw  (j�^  ]rw  (j�^  ]rw  (j�^  ]rw  (h	h�e]rw  (hh�e]rw  (hhe]rw  (j�^  ]rw  (h	he]rw  (hh�e]rw  (hhe]rw  (j�s  ]rw  (h	h�e]rw  (hh�eeee]r w  (hhee]r!w  (h!]r"w  (h#h$e]r#w  (h	he]r$w  (hh�e]r%w  (h)heeejw  jw  jw  jw  jw  jw  jw  jw  jw  ]r&w  (j�^  ]r'w  (j�^  ]r(w  (j�^  ]r)w  (h	h�e]r*w  (hh�e]r+w  (hhe]r,w  (j�^  ]r-w  (h	he]r.w  (hh�e]r/w  (hhe]r0w  (j�s  ]r1w  (h	h�e]r2w  (hh�eeee]r3w  (hhee]r4w  (h!]r5w  (h#h$e]r6w  (h	he]r7w  (hh�e]r8w  (h)heeej&w  j&w  j&w  j&w  ]r9w  (j�^  ]r:w  (j�^  ]r;w  (j�^  ]r<w  (h	h�e]r=w  (hh�e]r>w  (hhe]r?w  (j�^  ]r@w  (h	he]rAw  (hh�e]rBw  (hhe]rCw  (j�s  ]rDw  (h	h�e]rEw  (hh�eeee]rFw  (hhee]rGw  (h!]rHw  (h#h$e]rIw  (h	he]rJw  (hh�e]rKw  (h)heeej9w  ]rLw  (j�^  ]rMw  (j�^  ]rNw  (j�^  ]rOw  (h	h�e]rPw  (hh�e]rQw  (hhe]rRw  (j�^  ]rSw  (h	he]rTw  (hh�e]rUw  (hhe]rVw  (j�s  ]rWw  (h	h�e]rXw  (hh�eeee]rYw  (hhee]rZw  (h!]r[w  (h#h$e]r\w  (h	he]r]w  (hh�e]r^w  (h)heee]r_w  (j�^  ]r`w  (j�^  ]raw  (j�^  ]rbw  (h	h�e]rcw  (hh�e]rdw  (hhe]rew  (j�^  ]rfw  (h	he]rgw  (hh�e]rhw  (hhe]riw  (j�s  ]rjw  (h	h�e]rkw  (hh�eeee]rlw  (hhee]rmw  (h!]rnw  (h#h$e]row  (h	he]rpw  (hh�e]rqw  (h)heee]rrw  (j�^  ]rsw  (j�^  ]rtw  (j�^  ]ruw  (h	h�e]rvw  (hh�e]rww  (hhe]rxw  (j�^  ]ryw  (h	he]rzw  (hh�e]r{w  (hhe]r|w  (X	   Next-Mover}w  ]r~w  (h	h�e]rw  (hh�eeee]r�w  (hhee]r�w  (h!]r�w  (h#h$e]r�w  (h	he]r�w  (hh�e]r�w  (h)heee]r�w  (j�^  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (h	h�e]r�w  (hh�e]r�w  (hhe]r�w  (j�^  ]r�w  (h	he]r�w  (hh�e]r�w  (hhe]r�w  (j}w  ]r�w  (h	h�e]r�w  (hh�eeee]r�w  (hhee]r�w  (h!]r�w  (h#h$e]r�w  (h	he]r�w  (hh�e]r�w  (h)heeej�w  j�w  j�w  j�w  j�w  j�w  j�w  j�w  j�w  j�w  j�w  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (h	h�e]r�w  (hh�e]r�w  (hhe]r�w  (j�^  ]r�w  (h	he]r�w  (hh�e]r�w  (hhe]r�w  (j}w  ]r�w  (h	h�e]r�w  (hh�eeee]r�w  (hhee]r�w  (h!]r�w  (h#h$e]r�w  (h	he]r�w  (hh�e]r�w  (h)heeej�w  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (h	h�e]r�w  (hh�e]r�w  (hhe]r�w  (j�^  ]r�w  (h	he]r�w  (hh�e]r�w  (hhe]r�w  (j}w  ]r�w  (h	h�e]r�w  (hh�eeee]r�w  (hhee]r�w  (h!]r�w  (h#h$e]r�w  (h	he]r�w  (hh�e]r�w  (h)heeej�w  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (h	h�e]r�w  (hh�e]r�w  (hhe]r�w  (j�^  ]r�w  (h	he]r�w  (hh�e]r�w  (hhe]r�w  (j}w  ]r�w  (h	h�e]r�w  (hh�eeee]r�w  (hhee]r�w  (h!]r�w  (h#h$e]r�w  (h	he]r�w  (hh�e]r�w  (h)heeej�w  j�w  j�w  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (h	h�e]r�w  (hh�e]r�w  (hhe]r�w  (j�^  ]r�w  (h	he]r�w  (hh�e]r�w  (hhe]r�w  (j}w  ]r�w  (h	h�e]r�w  (hh�eeee]r�w  (hhee]r�w  (h!]r�w  (h#h$e]r�w  (h	he]r�w  (hh�e]r�w  (h)heeej�w  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (h	h�e]r�w  (hh�e]r�w  (hhe]r�w  (j�^  ]r�w  (h	he]r�w  (hh�e]r�w  (hhe]r�w  (j}w  ]r�w  (h	h�e]r�w  (hh�eeee]r�w  (hhee]r�w  (h!]r�w  (h#h$e]r�w  (h	he]r�w  (hh�e]r�w  (h)heee]r�w  (j�^  ]r�w  (j�^  ]r�w  (j�^  ]r�w  (h	h�e]r�w  (hh�e]r�w  (hhe]r�w  (j�^  ]r�w  (h	he]r x  (hh�e]rx  (hhe]rx  (j}w  ]rx  (h	h�e]rx  (hh�eeee]rx  (hhee]rx  (h!]rx  (h#h$e]rx  (h	he]r	x  (hh�e]r
x  (h)heeej�w  j�w  j�w  j�w  ]rx  (j�^  ]rx  (j�^  ]rx  (j�^  ]rx  (h	h�e]rx  (hh�e]rx  (hhe]rx  (j�^  ]rx  (h	he]rx  (hh�e]rx  (hhe]rx  (j}w  ]rx  (h	h�e]rx  (hh�eeee]rx  (hhee]rx  (h!]rx  (h#h$e]rx  (h	he]rx  (hh�e]rx  (h)heeejx  jx  jx  ]rx  (j�^  ]rx  (j�^  ]r x  (j�^  ]r!x  (h	h�e]r"x  (hh�e]r#x  (hhe]r$x  (j�^  ]r%x  (h	he]r&x  (hh�e]r'x  (hhe]r(x  (j}w  ]r)x  (h	h�e]r*x  (hh�eeee]r+x  (hhee]r,x  (h!]r-x  (h#h$e]r.x  (h	he]r/x  (hh�e]r0x  (h)heeejx  jx  jx  jx  jx  jx  ]r1x  (j�^  ]r2x  (j�^  ]r3x  (j�^  ]r4x  (h	h�e]r5x  (hh�e]r6x  (hhe]r7x  (j�^  ]r8x  (h	he]r9x  (hh�e]r:x  (hhe]r;x  (j}w  ]r<x  (h	h�e]r=x  (hh�eeee]r>x  (hhee]r?x  (h!]r@x  (h#h$e]rAx  (h	he]rBx  (hh�e]rCx  (h)heeej1x  j1x  j1x  ]rDx  (j�^  ]rEx  (j�^  ]rFx  (j�^  ]rGx  (h	h�e]rHx  (hh�e]rIx  (hhe]rJx  (j�^  ]rKx  (h	he]rLx  (hh�e]rMx  (hhe]rNx  (j}w  ]rOx  (h	h�e]rPx  (hh�eeee]rQx  (hhee]rRx  (h!]rSx  (h#h$e]rTx  (h	he]rUx  (hh�e]rVx  (h)heee]rWx  (j�^  ]rXx  (j�^  ]rYx  (j�^  ]rZx  (h	h�e]r[x  (hh�e]r\x  (hhe]r]x  (j�^  ]r^x  (h	he]r_x  (hh�e]r`x  (hhe]rax  (j}w  ]rbx  (h	h�e]rcx  (hh�eeee]rdx  (hhee]rex  (h!]rfx  (h#h$e]rgx  (h	he]rhx  (hh�e]rix  (h)heeejWx  jWx  ]rjx  (j�^  ]rkx  (j�^  ]rlx  (j�^  ]rmx  (h	h�e]rnx  (hh�e]rox  (hhe]rpx  (j�^  ]rqx  (h	he]rrx  (hh�e]rsx  (hhe]rtx  (j}w  ]rux  (h	h�e]rvx  (hh�eeee]rwx  (hhee]rxx  (h!]ryx  (h#h$e]rzx  (h	he]r{x  (hh�e]r|x  (h)heeejjx  ]r}x  (j�^  ]r~x  (j�^  ]rx  (j�^  ]r�x  (h	h�e]r�x  (hh�e]r�x  (hhe]r�x  (j�^  ]r�x  (h	he]r�x  (hh�e]r�x  (hhe]r�x  (j}w  ]r�x  (h	h�e]r�x  (hh�eeee]r�x  (hhee]r�x  (h!]r�x  (h#h$e]r�x  (h	he]r�x  (hh�e]r�x  (h)heeej}x  j}x  j}x  j}x  j}x  j}x  j}x  j}x  ]r�x  (j�^  ]r�x  (j�^  ]r�x  (j�^  ]r�x  (h	h�e]r�x  (hh�e]r�x  (hhe]r�x  (j�^  ]r�x  (h	he]r�x  (hh�e]r�x  (hhe]r�x  (j}w  ]r�x  (h	h�e]r�x  (hh�eeee]r�x  (hhee]r�x  (h!]r�x  (h#h$e]r�x  (h	he]r�x  (hh�e]r�x  (h)heeej�x  ]r�x  (j�^  ]r�x  (j�^  ]r�x  (j�^  ]r�x  (h	h�e]r�x  (hh�e]r�x  (hhe]r�x  (j�^  ]r�x  (h	he]r�x  (hh�e]r�x  (hhe]r�x  (j}w  ]r�x  (h	h�e]r�x  (hh�eeee]r�x  (hhee]r�x  (h!]r�x  (h#h$e]r�x  (h	he]r�x  (hh�e]r�x  (h)heee]r�x  (j�^  ]r�x  (j�^  ]r�x  (j�^  ]r�x  (h	h�e]r�x  (hh�e]r�x  (hhe]r�x  (j�^  ]r�x  (h	he]r�x  (hh�e]r�x  (hhe]r�x  (j}w  ]r�x  (h	h�e]r�x  (hh�eeee]r�x  (hhee]r�x  (h!]r�x  (h#h$e]r�x  (h	he]r�x  (hh�e]r�x  (h)heeej�x  j�x  ]r�x  (j�^  ]r�x  (j�^  ]r�x  (j�^  ]r�x  (h	h�e]r�x  (hh�e]r�x  (hhe]r�x  (j�^  ]r�x  (h	he]r�x  (hh�e]r�x  (hhe]r�x  (j}w  ]r�x  (h	h�e]r�x  (hh�eeee]r�x  (hhee]r�x  (h!]r�x  (h#h$e]r�x  (h	he]r�x  (hh�e]r�x  (h)heeej�x  j�x  ]r�x  (j�^  ]r�x  (j�^  ]r�x  (j�^  ]r�x  (h	h�e]r�x  (hh�e]r�x  (hhe]r�x  (j�^  ]r�x  (h	he]r�x  (hh�e]r�x  (hhe]r�x  (j}w  ]r�x  (h	h�e]r�x  (hh�eeee]r�x  (hhee]r�x  (h!]r�x  (h#h$e]r�x  (h	he]r�x  (hh�e]r�x  (h)heeej�x  ]r�x  (j�^  ]r�x  (j�^  ]r�x  (j�^  ]r�x  (h	h�e]r�x  (hh�e]r�x  (hhe]r�x  (j�^  ]r�x  (h	he]r�x  (hh�e]r�x  (hhe]r�x  (j}w  ]r�x  (h	h�e]r�x  (hh�eeee]r�x  (hhee]r�x  (h!]r�x  (h#h$e]r�x  (h	he]r y  (hh�e]ry  (h)heeej�x  j�x  j�x  j�x  ]ry  (j�^  ]ry  (j�^  ]ry  (j�^  ]ry  (h	h�e]ry  (hh�e]ry  (hhe]ry  (j�^  ]r	y  (h	he]r
y  (hh�e]ry  (hhe]ry  (j}w  ]ry  (h	h�e]ry  (hh�eeee]ry  (hhee]ry  (h!]ry  (h#h$e]ry  (h	he]ry  (hh�e]ry  (h)heeejy  jy  jy  jy  jy  jy  jy  jy  jy  ]ry  (j�^  ]ry  (j�^  ]ry  (j�^  ]ry  (h	h�e]ry  (hh�e]ry  (hhe]ry  (j�^  ]ry  (h	he]ry  (hh�e]ry  (hhe]ry  (j}w  ]r y  (h	h�e]r!y  (hh�eeee]r"y  (hhee]r#y  (h!]r$y  (h#h$e]r%y  (h	he]r&y  (hh�e]r'y  (h)heeejy  jy  jy  jy  jy  jy  jy  jy  ]r(y  (j�^  ]r)y  (j�^  ]r*y  (j�^  ]r+y  (h	h�e]r,y  (hh�e]r-y  (hhe]r.y  (j�^  ]r/y  (h	he]r0y  (hh�e]r1y  (hhe]r2y  (j}w  ]r3y  (h	h�e]r4y  (hh�eeee]r5y  (hhee]r6y  (h!]r7y  (h#h$e]r8y  (h	he]r9y  (hh�e]r:y  (h)heee]r;y  (j�^  ]r<y  (j�^  ]r=y  (j�^  ]r>y  (h	h�e]r?y  (hh�e]r@y  (hhe]rAy  (j�^  ]rBy  (h	he]rCy  (hh�e]rDy  (hhe]rEy  (j}w  ]rFy  (h	h�e]rGy  (hh�eeee]rHy  (hhee]rIy  (h!]rJy  (h#h$e]rKy  (h	he]rLy  (hh�e]rMy  (h)heeej;y  j;y  j;y  j;y  j;y  j;y  j;y  j;y  ]rNy  (j�^  ]rOy  (j�^  ]rPy  (j�^  ]rQy  (h	h�e]rRy  (hh�e]rSy  (hhe]rTy  (j�^  ]rUy  (h	he]rVy  (hh�e]rWy  (hhe]rXy  (j}w  ]rYy  (h	h�e]rZy  (hh�eeee]r[y  (hhee]r\y  (h!]r]y  (h#h$e]r^y  (h	he]r_y  (hh�e]r`y  (h)heeejNy  jNy  jNy  jNy  jNy  jNy  jNy  jNy  ]ray  (j�^  ]rby  (j�^  ]rcy  (j�^  ]rdy  (h	h�e]rey  (hh�e]rfy  (hhe]rgy  (j�^  ]rhy  (h	he]riy  (hh�e]rjy  (hhe]rky  (j}w  ]rly  (h	h�e]rmy  (hh�eeee]rny  (hhee]roy  (h!]rpy  (h#h$e]rqy  (h	he]rry  (hh�e]rsy  (h)heeejay  jay  jay  jay  jay  jay  ]rty  (j�^  ]ruy  (j�^  ]rvy  (j�^  ]rwy  (h	h�e]rxy  (hh�e]ryy  (hhe]rzy  (j�^  ]r{y  (h	he]r|y  (hh�e]r}y  (hhe]r~y  (j}w  ]ry  (h	h�e]r�y  (hh�eeee]r�y  (hhee]r�y  (h!]r�y  (h#h$e]r�y  (h	he]r�y  (hh�e]r�y  (h)heee]r�y  (j�^  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (h	h�e]r�y  (hh�e]r�y  (hhe]r�y  (j�^  ]r�y  (h	he]r�y  (hh�e]r�y  (hhe]r�y  (j}w  ]r�y  (h	h�e]r�y  (hh�eeee]r�y  (hhee]r�y  (h!]r�y  (h#h$e]r�y  (h	he]r�y  (hh�e]r�y  (h)heee]r�y  (j�^  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (h	h�e]r�y  (hh�e]r�y  (hhe]r�y  (j�^  ]r�y  (h	he]r�y  (hh�e]r�y  (hhe]r�y  (j}w  ]r�y  (h	h�e]r�y  (hh�eeee]r�y  (hhee]r�y  (h!]r�y  (h#h$e]r�y  (h	he]r�y  (hh�e]r�y  (h)heeej�y  j�y  j�y  j�y  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (h	h�e]r�y  (hh�e]r�y  (hhe]r�y  (j�^  ]r�y  (h	he]r�y  (hh�e]r�y  (hhe]r�y  (j}w  ]r�y  (h	h�e]r�y  (hh�eeee]r�y  (hhee]r�y  (h!]r�y  (h#h$e]r�y  (h	he]r�y  (hh�e]r�y  (h)heeej�y  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (h	h�e]r�y  (hh�e]r�y  (hhe]r�y  (j�^  ]r�y  (h	he]r�y  (hh�e]r�y  (hhe]r�y  (j}w  ]r�y  (h	h�e]r�y  (hh�eeee]r�y  (hhee]r�y  (h!]r�y  (h#h$e]r�y  (h	he]r�y  (hh�e]r�y  (h)heeej�y  j�y  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (h	h�e]r�y  (hh�e]r�y  (hhe]r�y  (j�^  ]r�y  (h	he]r�y  (hh�e]r�y  (hhe]r�y  (j}w  ]r�y  (h	h�e]r�y  (hh�eeee]r�y  (hhee]r�y  (h!]r�y  (h#h$e]r�y  (h	he]r�y  (hh�e]r�y  (h)heeej�y  j�y  j�y  j�y  j�y  j�y  j�y  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (h	h�e]r�y  (hh�e]r�y  (hhe]r�y  (j�^  ]r�y  (h	he]r�y  (hh�e]r�y  (hhe]r�y  (j}w  ]r�y  (h	h�e]r�y  (hh�eeee]r�y  (hhee]r�y  (h!]r�y  (h#h$e]r�y  (h	he]r�y  (hh�e]r�y  (h)heeej�y  j�y  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (j�^  ]r�y  (h	h�e]r�y  (hh�e]r�y  (hhe]r�y  (j�^  ]r z  (h	he]rz  (hh�e]rz  (hhe]rz  (j}w  ]rz  (h	h�e]rz  (hh�eeee]rz  (hhee]rz  (h!]rz  (h#h$e]r	z  (h	he]r
z  (hh�e]rz  (h)heeej�y  j�y  j�y  ]rz  (j�^  ]rz  (j�^  ]rz  (j�^  ]rz  (h	h�e]rz  (hh�e]rz  (hhe]rz  (j�^  ]rz  (h	he]rz  (hh�e]rz  (hhe]rz  (j}w  ]rz  (h	h�e]rz  (hh�eeee]rz  (hhee]rz  (h!]rz  (h#h$e]rz  (h	he]rz  (hh�e]rz  (h)heeejz  jz  ]rz  (j�^  ]r z  (j�^  ]r!z  (j�^  ]r"z  (h	h�e]r#z  (hh�e]r$z  (hhe]r%z  (j�^  ]r&z  (h	he]r'z  (hh�e]r(z  (hhe]r)z  (j}w  ]r*z  (h	h�e]r+z  (hh�eeee]r,z  (hhee]r-z  (h!]r.z  (h#h$e]r/z  (h	he]r0z  (hh�e]r1z  (h)heeejz  jz  ]r2z  (j�^  ]r3z  (j�^  ]r4z  (j�^  ]r5z  (h	h�e]r6z  (hh�e]r7z  (hhe]r8z  (j�^  ]r9z  (h	he]r:z  (hh�e]r;z  (hhe]r<z  (j}w  ]r=z  (h	h�e]r>z  (hh�eeee]r?z  (hhee]r@z  (h!]rAz  (h#h$e]rBz  (h	he]rCz  (hh�e]rDz  (h)heeej2z  j2z  ]rEz  (j�^  ]rFz  (j�^  ]rGz  (j�^  ]rHz  (h	h�e]rIz  (hh�e]rJz  (hhe]rKz  (j�^  ]rLz  (h	he]rMz  (hh�e]rNz  (hhe]rOz  (j}w  ]rPz  (h	h�e]rQz  (hh�eeee]rRz  (hhee]rSz  (h!]rTz  (h#h$e]rUz  (h	he]rVz  (hh�e]rWz  (h)heeejEz  ]rXz  (j�^  ]rYz  (j�^  ]rZz  (j�^  ]r[z  (h	h�e]r\z  (hh�e]r]z  (hhe]r^z  (j�^  ]r_z  (h	he]r`z  (hh�e]raz  (hhe]rbz  (j}w  ]rcz  (h	h�e]rdz  (hh�eeee]rez  (hhee]rfz  (h!]rgz  (h#h$e]rhz  (h	he]riz  (hh�e]rjz  (h)heeejXz  jXz  jXz  ]rkz  (j�^  ]rlz  (j�^  ]rmz  (j�^  ]rnz  (h	h�e]roz  (hh�e]rpz  (hhe]rqz  (j�^  ]rrz  (h	he]rsz  (hh�e]rtz  (hhe]ruz  (j}w  ]rvz  (h	h�e]rwz  (hh�eeee]rxz  (hhee]ryz  (h!]rzz  (h#h$e]r{z  (h	he]r|z  (hh�e]r}z  (h)heeejkz  jkz  jkz  ]r~z  (j�^  ]rz  (j�^  ]r�z  (j�^  ]r�z  (h	h�e]r�z  (hh�e]r�z  (hhe]r�z  (j�^  ]r�z  (h	he]r�z  (hh�e]r�z  (hhe]r�z  (j}w  ]r�z  (h	h�e]r�z  (hh�eeee]r�z  (hhee]r�z  (h!]r�z  (h#h$e]r�z  (h	he]r�z  (hh�e]r�z  (h)heeej~z  j~z  j~z  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (h	h�e]r�z  (hh�e]r�z  (hhe]r�z  (j�^  ]r�z  (h	he]r�z  (hh�e]r�z  (hhe]r�z  (j}w  ]r�z  (h	h�e]r�z  (hh�eeee]r�z  (hhee]r�z  (h!]r�z  (h#h$e]r�z  (h	he]r�z  (hh�e]r�z  (h)heeej�z  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (h	h�e]r�z  (hh�e]r�z  (hhe]r�z  (j�^  ]r�z  (h	he]r�z  (hh�e]r�z  (hhe]r�z  (j}w  ]r�z  (h	h�e]r�z  (hh�eeee]r�z  (hhee]r�z  (h!]r�z  (h#h$e]r�z  (h	he]r�z  (hh�e]r�z  (h)heeej�z  j�z  j�z  j�z  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (h	h�e]r�z  (hh�e]r�z  (hhe]r�z  (j�^  ]r�z  (h	he]r�z  (hh�e]r�z  (hhe]r�z  (j}w  ]r�z  (h	h�e]r�z  (hh�eeee]r�z  (hhee]r�z  (h!]r�z  (h#h$e]r�z  (h	he]r�z  (hh�e]r�z  (h)heeej�z  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (h	h�e]r�z  (hh�e]r�z  (hhe]r�z  (j�^  ]r�z  (h	he]r�z  (hh�e]r�z  (hhe]r�z  (j}w  ]r�z  (h	h�e]r�z  (hh�eeee]r�z  (hhee]r�z  (h!]r�z  (h#h$e]r�z  (h	he]r�z  (hh�e]r�z  (h)heeej�z  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (h	h�e]r�z  (hh�e]r�z  (hhe]r�z  (j�^  ]r�z  (h	he]r�z  (hh�e]r�z  (hhe]r�z  (j}w  ]r�z  (h	h�e]r�z  (hh�eeee]r�z  (hhee]r�z  (h!]r�z  (h#h$e]r�z  (h	he]r�z  (hh�e]r�z  (h)heeej�z  j�z  j�z  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (j�^  ]r�z  (h	h�e]r�z  (hh�e]r�z  (hhe]r�z  (j�^  ]r�z  (h	h�e]r�z  (hh�e]r�z  (hhe]r�z  (j}w  ]r�z  (h	h�e]r�z  (hh�eeee]r�z  (hhee]r�z  (h!]r�z  (h#h$e]r {  (h	he]r{  (hh�e]r{  (h)heeej�z  ]r{  (j�^  ]r{  (j�^  ]r{  (j�^  ]r{  (h	h�e]r{  (hh�e]r{  (hhe]r	{  (j�^  ]r
{  (h	h�e]r{  (hh�e]r{  (hhe]r{  (j}w  ]r{  (h	h�e]r{  (hh�eeee]r{  (hhee]r{  (h!]r{  (h#h$e]r{  (h	he]r{  (hh�e]r{  (h)heeej{  j{  j{  ]r{  (j�^  ]r{  (j�^  ]r{  (j�^  ]r{  (h	h�e]r{  (hh�e]r{  (hhe]r{  (j�^  ]r{  (h	h�e]r{  (hh�e]r{  (hhe]r {  (j}w  ]r!{  (h	h�e]r"{  (hh�eeee]r#{  (hhee]r${  (h!]r%{  (h#h$e]r&{  (h	he]r'{  (hh�e]r({  (h)heeej{  j{  j{  j{  ]r){  (j�^  ]r*{  (j�^  ]r+{  (j�^  ]r,{  (h	h�e]r-{  (hh�e]r.{  (hhe]r/{  (j�^  ]r0{  (h	h�e]r1{  (hh�e]r2{  (hhe]r3{  (j}w  ]r4{  (h	h�e]r5{  (hh�eeee]r6{  (hhee]r7{  (h!]r8{  (h#h$e]r9{  (h	he]r:{  (hh�e]r;{  (h)heeej){  j){  ]r<{  (j�^  ]r={  (j�^  ]r>{  (j�^  ]r?{  (h	h�e]r@{  (hh�e]rA{  (hhe]rB{  (j�^  ]rC{  (h	h�e]rD{  (hh�e]rE{  (hhe]rF{  (j}w  ]rG{  (h	h�e]rH{  (hh�eeee]rI{  (hhee]rJ{  (h!]rK{  (h#h$e]rL{  (h	he]rM{  (hh�e]rN{  (h)heee]rO{  (j�^  ]rP{  (j�^  ]rQ{  (j�^  ]rR{  (h	h�e]rS{  (hh�e]rT{  (hhe]rU{  (j�^  ]rV{  (h	h�e]rW{  (hh�e]rX{  (hhe]rY{  (j}w  ]rZ{  (h	h�e]r[{  (hh�eeee]r\{  (hhee]r]{  (h!]r^{  (h#h$e]r_{  (h	he]r`{  (hh�e]ra{  (h)heeejO{  jO{  jO{  jO{  ]rb{  (j�^  ]rc{  (j�^  ]rd{  (j�^  ]re{  (h	h�e]rf{  (hh�e]rg{  (hhe]rh{  (j�^  ]ri{  (h	h�e]rj{  (hh�e]rk{  (hhe]rl{  (j}w  ]rm{  (h	h�e]rn{  (hh�eeee]ro{  (hhee]rp{  (h!]rq{  (h#h$e]rr{  (h	he]rs{  (hh�e]rt{  (h)heeejb{  ]ru{  (j�^  ]rv{  (j�^  ]rw{  (j�^  ]rx{  (h	h�e]ry{  (hh�e]rz{  (hhe]r{{  (j�^  ]r|{  (h	he]r}{  (hh�e]r~{  (hhe]r{  (j}w  ]r�{  (h	h�e]r�{  (hh�eeee]r�{  (hhee]r�{  (h!]r�{  (h#h$e]r�{  (h	he]r�{  (hh�e]r�{  (h)heeeju{  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (h	h�e]r�{  (hh�e]r�{  (hhe]r�{  (j�^  ]r�{  (h	he]r�{  (hh�e]r�{  (hhe]r�{  (j}w  ]r�{  (h	h�e]r�{  (hh�eeee]r�{  (hhee]r�{  (h!]r�{  (h#h$e]r�{  (h	he]r�{  (hh�e]r�{  (h)heeej�{  j�{  j�{  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (h	h�e]r�{  (hh�e]r�{  (hhe]r�{  (j�^  ]r�{  (h	he]r�{  (hh�e]r�{  (hhe]r�{  (j}w  ]r�{  (h	h�e]r�{  (hh�eeee]r�{  (hhee]r�{  (h!]r�{  (h#h$e]r�{  (h	he]r�{  (hh�e]r�{  (h)heeej�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (h	h�e]r�{  (hh�e]r�{  (hhe]r�{  (j�^  ]r�{  (h	he]r�{  (hh�e]r�{  (hhe]r�{  (j}w  ]r�{  (h	h�e]r�{  (hh�eeee]r�{  (hhee]r�{  (h!]r�{  (h#h$e]r�{  (h	he]r�{  (hh�e]r�{  (h)heee]r�{  (j�^  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (h	h�e]r�{  (hh�e]r�{  (hhe]r�{  (j�^  ]r�{  (h	he]r�{  (hh�e]r�{  (hhe]r�{  (j}w  ]r�{  (h	h�e]r�{  (hh�eeee]r�{  (hhee]r�{  (h!]r�{  (h#h$e]r�{  (h	he]r�{  (hh�e]r�{  (h)heee]r�{  (j�^  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (h	h�e]r�{  (hh�e]r�{  (hhe]r�{  (j�^  ]r�{  (h	he]r�{  (hh�e]r�{  (hhe]r�{  (j}w  ]r�{  (h	h�e]r�{  (hh�eeee]r�{  (hhee]r�{  (h!]r�{  (h#h$e]r�{  (h	he]r�{  (hh�e]r�{  (h)heeej�{  j�{  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (h	h�e]r�{  (hh�e]r�{  (hhe]r�{  (j�^  ]r�{  (h	he]r�{  (hh�e]r�{  (hhe]r�{  (j}w  ]r�{  (h	h�e]r�{  (hh�eeee]r�{  (hhee]r�{  (h!]r�{  (h#h$e]r�{  (h	he]r�{  (hh�e]r�{  (h)heeej�{  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (j�^  ]r�{  (h	h�e]r�{  (hh�e]r�{  (hhe]r |  (j�^  ]r|  (h	he]r|  (hh�e]r|  (hhe]r|  (j}w  ]r|  (h	h�e]r|  (hh�eeee]r|  (hhee]r|  (h!]r	|  (h#h$e]r
|  (h	he]r|  (hh�e]r|  (h)heeej�{  ]r|  (j�^  ]r|  (j�^  ]r|  (j�^  ]r|  (h	h�e]r|  (hh�e]r|  (hhe]r|  (j�^  ]r|  (h	he]r|  (hh�e]r|  (hhe]r|  (j}w  ]r|  (h	h�e]r|  (hh�eeee]r|  (hhee]r|  (h!]r|  (h#h$e]r|  (h	he]r|  (hh�e]r|  (h)heeej|  j|  ]r |  (j�^  ]r!|  (j�^  ]r"|  (j�^  ]r#|  (h	h�e]r$|  (hh�e]r%|  (hhe]r&|  (j�^  ]r'|  (h	he]r(|  (hh�e]r)|  (hhe]r*|  (j}w  ]r+|  (h	h�e]r,|  (hh�eeee]r-|  (hhee]r.|  (h!]r/|  (h#h$e]r0|  (h	he]r1|  (hh�e]r2|  (h)heeej |  j |  j |  j |  j |  j |  ]r3|  (j�^  ]r4|  (j�^  ]r5|  (j�^  ]r6|  (h	h�e]r7|  (hh�e]r8|  (hhe]r9|  (j�^  ]r:|  (h	he]r;|  (hh�e]r<|  (hhe]r=|  (j}w  ]r>|  (h	h�e]r?|  (hh�eeee]r@|  (hhee]rA|  (h!]rB|  (h#h$e]rC|  (h	he]rD|  (hh�e]rE|  (h)heeej3|  j3|  ]rF|  (j�^  ]rG|  (j�^  ]rH|  (j�^  ]rI|  (h	h�e]rJ|  (hh�e]rK|  (hhe]rL|  (j�^  ]rM|  (h	he]rN|  (hh�e]rO|  (hhe]rP|  (j}w  ]rQ|  (h	h�e]rR|  (hh�eeee]rS|  (hhee]rT|  (h!]rU|  (h#h$e]rV|  (h	he]rW|  (hh�e]rX|  (h)heee]rY|  (j�^  ]rZ|  (j�^  ]r[|  (j�^  ]r\|  (h	h�e]r]|  (hh�e]r^|  (hhe]r_|  (j�^  ]r`|  (h	he]ra|  (hh�e]rb|  (hhe]rc|  (j}w  ]rd|  (h	h�e]re|  (hh�eeee]rf|  (hhee]rg|  (h!]rh|  (h#h$e]ri|  (h	he]rj|  (hh�e]rk|  (h)heeejY|  jY|  jY|  jY|  jY|  ]rl|  (j�^  ]rm|  (j�^  ]rn|  (j�^  ]ro|  (h	h�e]rp|  (hh�e]rq|  (hhe]rr|  (j�^  ]rs|  (h	he]rt|  (hh�e]ru|  (hhe]rv|  (j}w  ]rw|  (h	h�e]rx|  (hh�eeee]ry|  (hhee]rz|  (h!]r{|  (h#h$e]r||  (h	he]r}|  (hh�e]r~|  (h)heee]r|  (j�^  ]r�|  (j�^  ]r�|  (j�^  ]r�|  (h	h�e]r�|  (hh�e]r�|  (hhe]r�|  (j�^  ]r�|  (h	he]r�|  (hh�e]r�|  (hhe]r�|  (j}w  ]r�|  (h	h�e]r�|  (hh�eeee]r�|  (hhee]r�|  (h!]r�|  (h#h$e]r�|  (h	he]r�|  (hh�e]r�|  (h)heee]r�|  (j�^  ]r�|  (j�^  ]r�|  (j�^  ]r�|  (h	h�e]r�|  (hh�e]r�|  (hhe]r�|  (j�^  ]r�|  (h	he]r�|  (hh�e]r�|  (hhe]r�|  (j}w  ]r�|  (h	h�e]r�|  (hh�eeee]r�|  (hhee]r�|  (h!]r�|  (h#h$e]r�|  (h	he]r�|  (hh�e]r�|  (h)heee]r�|  (j�^  ]r�|  (j�^  ]r�|  (j�^  ]r�|  (h	h�e]r�|  (hh�e]r�|  (hhe]r�|  (j�^  ]r�|  (h	he]r�|  (hh�e]r�|  (hhe]r�|  (j}w  ]r�|  (h	h�e]r�|  (hh�eeee]r�|  (hhee]r�|  (h!]r�|  (h#h$e]r�|  (h	he]r�|  (hh�e]r�|  (h)heeej�|  j�|  j�|  j�|  j�|  ]r�|  (j�^  ]r�|  (j�^  ]r�|  (j�^  ]r�|  (h	h�e]r�|  (hh�e]r�|  (hhe]r�|  (j�^  ]r�|  (h	he]r�|  (hh�e]r�|  (hhe]r�|  (j}w  ]r�|  (h	h�e]r�|  (hh�eeee]r�|  (hhee]r�|  (h!]r�|  (h#h$e]r�|  (h	he]r�|  (hh�e]r�|  (h)heeej�|  j�|  j�|  j�|  j�|  j�|  j�|  ]r�|  (j�^  ]r�|  (j�^  ]r�|  (j�^  ]r�|  (h	h�e]r�|  (hh�e]r�|  (hhe]r�|  (j�^  ]r�|  (h	he]r�|  (hh�e]r�|  (hhe]r�|  (j}w  ]r�|  (h	h�e]r�|  (hh�eeee]r�|  (hhee]r�|  (h!]r�|  (h#h$e]r�|  (h	he]r�|  (hh�e]r�|  (h)heeej�|  j�|  j�|  j�|  ]r�|  (j�^  ]r�|  (j�^  ]r�|  (j�^  ]r�|  (h	h�e]r�|  (hh�e]r�|  (hhe]r�|  (j�^  ]r�|  (h	he]r�|  (hh�e]r�|  (hhe]r�|  (j}w  ]r�|  (h	h�e]r�|  (hh�eeee]r�|  (hhee]r�|  (h!]r�|  (h#h$e]r�|  (h	he]r�|  (hh�e]r�|  (h)heeej�|  ]r�|  (j�^  ]r�|  (j�^  ]r�|  (j�^  ]r�|  (h	h�e]r�|  (hh�e]r�|  (hhe]r�|  (j�^  ]r�|  (h	he]r�|  (hh�e]r�|  (hhe]r�|  (j}w  ]r�|  (h	h�e]r�|  (hh�eeee]r�|  (hhee]r�|  (h!]r }  (h#h$e]r}  (h	he]r}  (hh�e]r}  (h)heeej�|  j�|  j�|  j�|  j�|  j�|  j�|  j�|  j�|  j�|  ]r}  (j�^  ]r}  (j�^  ]r}  (j�^  ]r}  (h	h�e]r}  (hh�e]r	}  (hhe]r
}  (j�^  ]r}  (h	he]r}  (hh�e]r}  (hhe]r}  (j}w  ]r}  (h	h�e]r}  (hh�eeee]r}  (hhee]r}  (h!]r}  (h#h$e]r}  (h	he]r}  (hh�e]r}  (h)heeej}  j}  j}  j}  j}  j}  j}  j}  j}  j}  ]r}  (j�^  ]r}  (j�^  ]r}  (j�^  ]r}  (h	h�e]r}  (hh�e]r}  (hhe]r}  (j�^  ]r}  (h	he]r}  (hh�e]r }  (hhe]r!}  (j}w  ]r"}  (h	h�e]r#}  (hh�eeee]r$}  (hhee]r%}  (h!]r&}  (h#h$e]r'}  (h	he]r(}  (hh�e]r)}  (h)heee]r*}  (j�^  ]r+}  (j�^  ]r,}  (j�^  ]r-}  (h	h�e]r.}  (hh�e]r/}  (hhe]r0}  (j�^  ]r1}  (h	he]r2}  (hh�e]r3}  (hhe]r4}  (j}w  ]r5}  (h	h�e]r6}  (hh�eeee]r7}  (hhee]r8}  (h!]r9}  (h#h$e]r:}  (h	he]r;}  (hh�e]r<}  (h)heeej*}  j*}  j*}  j*}  j*}  j*}  j*}  j*}  j*}  j*}  j*}  j*}  j*}  ]r=}  (j�^  ]r>}  (j�^  ]r?}  (j�^  ]r@}  (h	h�e]rA}  (hh�e]rB}  (hhe]rC}  (j�^  ]rD}  (h	he]rE}  (hh�e]rF}  (hhe]rG}  (j}w  ]rH}  (h	h�e]rI}  (hh�eeee]rJ}  (hhee]rK}  (h!]rL}  (h#h$e]rM}  (h	he]rN}  (hh�e]rO}  (h)heee]rP}  (j�^  ]rQ}  (j�^  ]rR}  (j�^  ]rS}  (h	h�e]rT}  (hh�e]rU}  (hhe]rV}  (j�^  ]rW}  (h	he]rX}  (hh�e]rY}  (hhe]rZ}  (j}w  ]r[}  (h	h�e]r\}  (hh�eeee]r]}  (hhee]r^}  (h!]r_}  (h#h$e]r`}  (h	he]ra}  (hh�e]rb}  (h)heee]rc}  (j�^  ]rd}  (j�^  ]re}  (j�^  ]rf}  (h	h�e]rg}  (hh�e]rh}  (hhe]ri}  (j�^  ]rj}  (h	he]rk}  (hh�e]rl}  (hhe]rm}  (j}w  ]rn}  (h	h�e]ro}  (hh�eeee]rp}  (hhee]rq}  (h!]rr}  (h#h$e]rs}  (h	he]rt}  (hh�e]ru}  (h)heeejc}  ]rv}  (j�^  ]rw}  (j�^  ]rx}  (j�^  ]ry}  (h	h�e]rz}  (hh�e]r{}  (hhe]r|}  (j�^  ]r}}  (h	he]r~}  (hh�e]r}  (hhe]r�}  (j}w  ]r�}  (h	h�e]r�}  (hh�eeee]r�}  (hhee]r�}  (h!]r�}  (h#h$e]r�}  (h	he]r�}  (hh�e]r�}  (h)heee]r�}  (j�^  ]r�}  (j�^  ]r�}  (j�^  ]r�}  (h	h�e]r�}  (hh�e]r�}  (hhe]r�}  (j�^  ]r�}  (h	he]r�}  (hh�e]r�}  (hhe]r�}  (j}w  ]r�}  (h	h�e]r�}  (hh�eeee]r�}  (hhee]r�}  (h!]r�}  (h#h$e]r�}  (h	he]r�}  (hh�e]r�}  (h)heee]r�}  (j�^  ]r�}  (j�^  ]r�}  (j�^  ]r�}  (h	h�e]r�}  (hh�e]r�}  (hhe]r�}  (j�^  ]r�}  (h	he]r�}  (hh�e]r�}  (hhe]r�}  (j}w  ]r�}  (h	h�e]r�}  (hh�eeee]r�}  (hhee]r�}  (h!]r�}  (h#h$e]r�}  (h	he]r�}  (hh�e]r�}  (h)heeej�}  ]r�}  (j�^  ]r�}  (j�^  ]r�}  (j�^  ]r�}  (h	h�e]r�}  (hh�e]r�}  (hhe]r�}  (j�^  ]r�}  (h	h�e]r�}  (hh�e]r�}  (hhe]r�}  (j}w  ]r�}  (h	h�e]r�}  (hh�eeee]r�}  (hhee]r�}  (h!]r�}  (h#h$e]r�}  (h	he]r�}  (hh�e]r�}  (h)heee]r�}  (j�^  ]r�}  (j�^  ]r�}  (j�^  ]r�}  (h	h�e]r�}  (hh�e]r�}  (hhe]r�}  (j�^  ]r�}  (h	h�e]r�}  (hh�e]r�}  (hhe]r�}  (j}w  ]r�}  (h	h�e]r�}  (hh�eeee]r�}  (hhee]r�}  (h!]r�}  (h#h$e]r�}  (h	he]r�}  (hh�e]r�}  (h)heeej�}  j�}  j�}  j�}  ]r�}  (j�^  ]r�}  (j�^  ]r�}  (j�^  ]r�}  (h	h�e]r�}  (hh�e]r�}  (hhe]r�}  (j�^  ]r�}  (h	h�e]r�}  (hh�e]r�}  (hhe]r�}  (j}w  ]r�}  (h	h�e]r�}  (hh�eeee]r�}  (hhee]r�}  (h!]r�}  (h#h$e]r�}  (h	he]r�}  (hh�e]r�}  (h)heee]r�}  (j�^  ]r�}  (j�^  ]r�}  (j�^  ]r�}  (h	h�e]r�}  (hh�e]r�}  (hhe]r�}  (j�^  ]r�}  (h	h�e]r�}  (hh�e]r�}  (hhe]r�}  (j}w  ]r�}  (h	h�e]r�}  (hh�eeee]r�}  (hhee]r�}  (h!]r�}  (h#h$e]r�}  (h	he]r�}  (hh�e]r�}  (h)heeej�}  ]r�}  (j�^  ]r�}  (j�^  ]r�}  (j�^  ]r�}  (h	h�e]r�}  (hh�e]r ~  (hhe]r~  (j�^  ]r~  (h	h�e]r~  (hh�e]r~  (hhe]r~  (j}w  ]r~  (h	h�e]r~  (hh�eeee]r~  (hhee]r	~  (h!]r
~  (h#h$e]r~  (h	he]r~  (hh�e]r~  (h)heeej�}  ]r~  (j�^  ]r~  (j�^  ]r~  (j�^  ]r~  (h	h�e]r~  (hh�e]r~  (hhe]r~  (j�^  ]r~  (h	h�e]r~  (hh�e]r~  (hhe]r~  (j}w  ]r~  (h	h�e]r~  (hh�eeee]r~  (hhee]r~  (h!]r~  (h#h$e]r~  (h	he]r~  (hh�e]r ~  (h)heeej~  j~  j~  ]r!~  (j�^  ]r"~  (j�^  ]r#~  (j�^  ]r$~  (h	h�e]r%~  (hh�e]r&~  (hhe]r'~  (j�^  ]r(~  (h	h�e]r)~  (hh�e]r*~  (hhe]r+~  (j}w  ]r,~  (h	h�e]r-~  (hh�eeee]r.~  (hhee]r/~  (h!]r0~  (h#h$e]r1~  (h	he]r2~  (hh�e]r3~  (h)heeej!~  j!~  j!~  j!~  j!~  j!~  ]r4~  (j�^  ]r5~  (j�^  ]r6~  (j�^  ]r7~  (h	h�e]r8~  (hh�e]r9~  (hhe]r:~  (j�^  ]r;~  (h	h�e]r<~  (hh�e]r=~  (hhe]r>~  (j}w  ]r?~  (h	h�e]r@~  (hh�eeee]rA~  (hhee]rB~  (h!]rC~  (h#h$e]rD~  (h	he]rE~  (hh�e]rF~  (h)heeej4~  j4~  ]rG~  (j�^  ]rH~  (j�^  ]rI~  (j�^  ]rJ~  (h	h�e]rK~  (hh�e]rL~  (hhe]rM~  (j�^  ]rN~  (h	h�e]rO~  (hh�e]rP~  (hhe]rQ~  (j}w  ]rR~  (h	h�e]rS~  (hh�eeee]rT~  (hhee]rU~  (h!]rV~  (h#h$e]rW~  (h	he]rX~  (hh�e]rY~  (h)heeejG~  jG~  ]rZ~  (j�^  ]r[~  (j�^  ]r\~  (j�^  ]r]~  (h	h�e]r^~  (hh�e]r_~  (hhe]r`~  (j�^  ]ra~  (h	h�e]rb~  (hh�e]rc~  (hhe]rd~  (j}w  ]re~  (h	h�e]rf~  (hh�eeee]rg~  (hhee]rh~  (h!]ri~  (h#h$e]rj~  (h	he]rk~  (hh�e]rl~  (h)heeejZ~  ]rm~  (j�^  ]rn~  (j�^  ]ro~  (j�^  ]rp~  (h	h�e]rq~  (hh�e]rr~  (hhe]rs~  (j�^  ]rt~  (h	h�e]ru~  (hh�e]rv~  (hhe]rw~  (j}w  ]rx~  (h	h�e]ry~  (hh�eeee]rz~  (hhee]r{~  (h!]r|~  (h#h$e]r}~  (h	he]r~~  (hh�e]r~  (h)heeejm~  jm~  jm~  jm~  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j}w  ]r�~  (h	h�e]r�~  (hh�eeee]r�~  (hhee]r�~  (h!]r�~  (h#h$e]r�~  (h	he]r�~  (hh�e]r�~  (h)heee]r�~  (j�^  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j}w  ]r�~  (h	h�e]r�~  (hh�eeee]r�~  (hhee]r�~  (h!]r�~  (h#h$e]r�~  (h	he]r�~  (hh�e]r�~  (h)heeej�~  j�~  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j}w  ]r�~  (h	h�e]r�~  (hh�eeee]r�~  (hhee]r�~  (h!]r�~  (h#h$e]r�~  (h	he]r�~  (hh�e]r�~  (h)heeej�~  j�~  j�~  j�~  j�~  j�~  j�~  j�~  j�~  j�~  j�~  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j}w  ]r�~  (h	h�e]r�~  (hh�eeee]r�~  (hhee]r�~  (h!]r�~  (h#h$e]r�~  (h	he]r�~  (hh�e]r�~  (h)heeej�~  j�~  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j}w  ]r�~  (h	h�e]r�~  (hh�eeee]r�~  (hhee]r�~  (h!]r�~  (h#h$e]r�~  (h	he]r�~  (hh�e]r�~  (h)heeej�~  j�~  j�~  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j}w  ]r�~  (h	h�e]r�~  (hh�eeee]r�~  (hhee]r�~  (h!]r�~  (h#h$e]r�~  (h	he]r�~  (hh�e]r�~  (h)heeej�~  j�~  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j�^  ]r�~  (h	h�e]r�~  (hh�e]r�~  (hhe]r�~  (j}w  ]r�~  (h	h�e]r�~  (hh�eeee]r�~  (hhee]r   (h!]r  (h#h$e]r  (h	he]r  (hh�e]r  (h)heeej�~  j�~  j�~  j�~  ]r  (j�^  ]r  (j�^  ]r  (j�^  ]r  (h	h�e]r	  (hh�e]r
  (hhe]r  (j�^  ]r  (h	h�e]r  (hh�e]r  (hhe]r  (j}w  ]r  (h	h�e]r  (hh�eeee]r  (hhee]r  (h!]r  (h#h$e]r  (h	he]r  (hh�e]r  (h)heeej  j  ]r  (j�^  ]r  (j�^  ]r  (j�^  ]r  (h	h�e]r  (hh�e]r  (hhe]r  (j�^  ]r  (h	h�e]r   (hh�e]r!  (hhe]r"  (j}w  ]r#  (h	h�e]r$  (hh�eeee]r%  (hhee]r&  (h!]r'  (h#h$e]r(  (h	he]r)  (hh�e]r*  (h)heeej  j  j  j  j  j  j  j  ]r+  (j�^  ]r,  (j�^  ]r-  (j�^  ]r.  (h	h�e]r/  (hh�e]r0  (hhe]r1  (j�^  ]r2  (h	h�e]r3  (hh�e]r4  (hhe]r5  (j}w  ]r6  (h	h�e]r7  (hh�eeee]r8  (hhee]r9  (h!]r:  (h#h$e]r;  (h	he]r<  (hh�e]r=  (h)heeej+  ]r>  (j�^  ]r?  (j�^  ]r@  (j�^  ]rA  (h	h�e]rB  (hh�e]rC  (hhe]rD  (j�^  ]rE  (h	h�e]rF  (hh�e]rG  (hhe]rH  (j}w  ]rI  (h	h�e]rJ  (hh�eeee]rK  (hhee]rL  (h!]rM  (h#h$e]rN  (h	he]rO  (hh�e]rP  (h)heee]rQ  (j�^  ]rR  (j�^  ]rS  (j�^  ]rT  (h	h�e]rU  (hh�e]rV  (hhe]rW  (j�^  ]rX  (h	h�e]rY  (hh�e]rZ  (hhe]r[  (j}w  ]r\  (h	h�e]r]  (hh�eeee]r^  (hhee]r_  (h!]r`  (h#h$e]ra  (h	he]rb  (hh�e]rc  (h)heee]rd  (j�^  ]re  (j�^  ]rf  (j�^  ]rg  (h	h�e]rh  (hh�e]ri  (hhe]rj  (j�^  ]rk  (h	h�e]rl  (hh�e]rm  (hhe]rn  (j}w  ]ro  (h	h�e]rp  (hh�eeee]rq  (hhee]rr  (h!]rs  (h#h$e]rt  (h	he]ru  (hh�e]rv  (h)heee]rw  (j�^  ]rx  (j�^  ]ry  (j�^  ]rz  (h	h�e]r{  (hh�e]r|  (hhe]r}  (j�^  ]r~  (h	h�e]r  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej�  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r �  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r	�  (hhee]r
�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r �  (hh�e]r!�  (h)heeej�  j�  j�  j�  ]r"�  (j�^  ]r#�  (j�^  ]r$�  (j�^  ]r%�  (h	h�e]r&�  (hh�e]r'�  (hhe]r(�  (j�^  ]r)�  (h	h�e]r*�  (hh�e]r+�  (hhe]r,�  (j}w  ]r-�  (h	h�e]r.�  (hh�eeee]r/�  (hhee]r0�  (h!]r1�  (h#h$e]r2�  (h	he]r3�  (hh�e]r4�  (h)heee]r5�  (j�^  ]r6�  (j�^  ]r7�  (j�^  ]r8�  (h	h�e]r9�  (hh�e]r:�  (hhe]r;�  (j�^  ]r<�  (h	h�e]r=�  (hh�e]r>�  (hhe]r?�  (j}w  ]r@�  (h	h�e]rA�  (hh�eeee]rB�  (hhee]rC�  (h!]rD�  (h#h$e]rE�  (h	he]rF�  (hh�e]rG�  (h)heeej5�  ]rH�  (j�^  ]rI�  (j�^  ]rJ�  (j�^  ]rK�  (h	h�e]rL�  (hh�e]rM�  (hhe]rN�  (j�^  ]rO�  (h	h�e]rP�  (hh�e]rQ�  (hhe]rR�  (j}w  ]rS�  (h	h�e]rT�  (hh�eeee]rU�  (hhee]rV�  (h!]rW�  (h#h$e]rX�  (h	he]rY�  (hh�e]rZ�  (h)heeejH�  jH�  jH�  jH�  jH�  ]r[�  (j�^  ]r\�  (j�^  ]r]�  (j�^  ]r^�  (h	h�e]r_�  (hh�e]r`�  (hhe]ra�  (j�^  ]rb�  (h	h�e]rc�  (hh�e]rd�  (hhe]re�  (j}w  ]rf�  (h	h�e]rg�  (hh�eeee]rh�  (hhee]ri�  (h!]rj�  (h#h$e]rk�  (h	he]rl�  (hh�e]rm�  (h)heeej[�  j[�  j[�  ]rn�  (j�^  ]ro�  (j�^  ]rp�  (j�^  ]rq�  (h	h�e]rr�  (hh�e]rs�  (hhe]rt�  (j�^  ]ru�  (h	h�e]rv�  (hh�e]rw�  (hhe]rx�  (j}w  ]ry�  (h	h�e]rz�  (hh�eeee]r{�  (hhee]r|�  (h!]r}�  (h#h$e]r~�  (h	he]r�  (hh�e]r��  (h)heeejn�  jn�  jn�  jn�  jn�  jn�  jn�  jn�  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heee]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heee]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	h�e]r  (hh�e]rÀ  (hhe]rĀ  (j}w  ]rŀ  (h	h�e]rƀ  (hh�eeee]rǀ  (hhee]rȀ  (h!]rɀ  (h#h$e]rʀ  (h	he]rˀ  (hh�e]r̀  (h)heeej��  ]r̀  (j�^  ]r΀  (j�^  ]rπ  (j�^  ]rЀ  (h	h�e]rр  (hh�e]rҀ  (hhe]rӀ  (j�^  ]rԀ  (h	he]rՀ  (hh�e]rր  (hhe]r׀  (j}w  ]r؀  (h	h�e]rـ  (hh�eeee]rڀ  (hhee]rۀ  (h!]r܀  (h#h$e]r݀  (h	he]rހ  (hh�e]r߀  (h)heeej̀  j̀  j̀  j̀  j̀  j̀  j̀  j̀  ]r��  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r��  (h	he]r�  (hh�e]r�  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  j��  ]r�  (j�^  ]r�  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r �  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r	�  (h	h�e]r
�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r �  (h	he]r!�  (hh�e]r"�  (hhe]r#�  (j}w  ]r$�  (h	h�e]r%�  (hh�eeee]r&�  (hhee]r'�  (h!]r(�  (h#h$e]r)�  (h	he]r*�  (hh�e]r+�  (h)heeej�  j�  j�  ]r,�  (j�^  ]r-�  (j�^  ]r.�  (j�^  ]r/�  (h	h�e]r0�  (hh�e]r1�  (hhe]r2�  (j�^  ]r3�  (h	he]r4�  (hh�e]r5�  (hhe]r6�  (j}w  ]r7�  (h	h�e]r8�  (hh�eeee]r9�  (hhee]r:�  (h!]r;�  (h#h$e]r<�  (h	he]r=�  (hh�e]r>�  (h)heeej,�  j,�  j,�  j,�  j,�  ]r?�  (j�^  ]r@�  (j�^  ]rA�  (j�^  ]rB�  (h	h�e]rC�  (hh�e]rD�  (hhe]rE�  (j�^  ]rF�  (h	he]rG�  (hh�e]rH�  (hhe]rI�  (j}w  ]rJ�  (h	h�e]rK�  (hh�eeee]rL�  (hhee]rM�  (h!]rN�  (h#h$e]rO�  (h	he]rP�  (hh�e]rQ�  (h)heeej?�  j?�  j?�  j?�  j?�  j?�  j?�  j?�  ]rR�  (j�^  ]rS�  (j�^  ]rT�  (j�^  ]rU�  (h	h�e]rV�  (hh�e]rW�  (hhe]rX�  (j�^  ]rY�  (h	he]rZ�  (hh�e]r[�  (hhe]r\�  (j}w  ]r]�  (h	h�e]r^�  (hh�eeee]r_�  (hhee]r`�  (h!]ra�  (h#h$e]rb�  (h	he]rc�  (hh�e]rd�  (h)heeejR�  jR�  jR�  jR�  jR�  ]re�  (j�^  ]rf�  (j�^  ]rg�  (j�^  ]rh�  (h	h�e]ri�  (hh�e]rj�  (hhe]rk�  (j�^  ]rl�  (h	he]rm�  (hh�e]rn�  (hhe]ro�  (j}w  ]rp�  (h	h�e]rq�  (hh�eeee]rr�  (hhee]rs�  (h!]rt�  (h#h$e]ru�  (h	he]rv�  (hh�e]rw�  (h)heeeje�  je�  je�  je�  je�  je�  je�  je�  je�  je�  ]rx�  (j�^  ]ry�  (j�^  ]rz�  (j�^  ]r{�  (h	h�e]r|�  (hh�e]r}�  (hhe]r~�  (j�^  ]r�  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeejx�  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heee]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heee]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r  (hh�e]rÁ  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  ]rā  (j�^  ]rŁ  (j�^  ]rƁ  (j�^  ]rǁ  (h	h�e]rȁ  (hh�e]rɁ  (hhe]rʁ  (j�^  ]rˁ  (h	he]ŕ  (hh�e]ŕ  (hhe]r΁  (j}w  ]rρ  (h	h�e]rЁ  (hh�eeee]rс  (hhee]rҁ  (h!]rӁ  (h#h$e]rԁ  (h	he]rՁ  (hh�e]rց  (h)heeejā  jā  jā  jā  jā  ]rׁ  (j�^  ]r؁  (j�^  ]rف  (j�^  ]rځ  (h	h�e]rہ  (hh�e]r܁  (hhe]r݁  (j�^  ]rށ  (h	he]r߁  (hh�e]r��  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeejׁ  jׁ  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r��  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heee]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r �  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r	�  (hh�eeee]r
�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r �  (h	he]r!�  (hh�e]r"�  (h)heee]r#�  (j�^  ]r$�  (j�^  ]r%�  (j�^  ]r&�  (h	h�e]r'�  (hh�e]r(�  (hhe]r)�  (j�^  ]r*�  (h	he]r+�  (hh�e]r,�  (hhe]r-�  (j}w  ]r.�  (h	h�e]r/�  (hh�eeee]r0�  (hhee]r1�  (h!]r2�  (h#h$e]r3�  (h	he]r4�  (hh�e]r5�  (h)heee]r6�  (j�^  ]r7�  (j�^  ]r8�  (j�^  ]r9�  (h	h�e]r:�  (hh�e]r;�  (hhe]r<�  (j�^  ]r=�  (h	he]r>�  (hh�e]r?�  (hhe]r@�  (j}w  ]rA�  (h	h�e]rB�  (hh�eeee]rC�  (hhee]rD�  (h!]rE�  (h#h$e]rF�  (h	he]rG�  (hh�e]rH�  (h)heeej6�  j6�  j6�  ]rI�  (j�^  ]rJ�  (j�^  ]rK�  (j�^  ]rL�  (h	h�e]rM�  (hh�e]rN�  (hhe]rO�  (j�^  ]rP�  (h	he]rQ�  (hh�e]rR�  (hhe]rS�  (j}w  ]rT�  (h	h�e]rU�  (hh�eeee]rV�  (hhee]rW�  (h!]rX�  (h#h$e]rY�  (h	he]rZ�  (hh�e]r[�  (h)heeejI�  jI�  jI�  jI�  jI�  jI�  ]r\�  (j�^  ]r]�  (j�^  ]r^�  (j�^  ]r_�  (h	h�e]r`�  (hh�e]ra�  (hhe]rb�  (j�^  ]rc�  (h	he]rd�  (hh�e]re�  (hhe]rf�  (j}w  ]rg�  (h	h�e]rh�  (hh�eeee]ri�  (hhee]rj�  (h!]rk�  (h#h$e]rl�  (h	he]rm�  (hh�e]rn�  (h)heee]ro�  (j�^  ]rp�  (j�^  ]rq�  (j�^  ]rr�  (h	h�e]rs�  (hh�e]rt�  (hhe]ru�  (j�^  ]rv�  (h	he]rw�  (hh�e]rx�  (hhe]ry�  (j}w  ]rz�  (h	h�e]r{�  (hh�eeee]r|�  (hhee]r}�  (h!]r~�  (h#h$e]r�  (h	he]r��  (hh�e]r��  (h)heeejo�  jo�  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heee]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r  (h	he]rÂ  (hh�e]rĂ  (hhe]rł  (j}w  ]rƂ  (h	h�e]rǂ  (hh�eeee]rȂ  (hhee]rɂ  (h!]rʂ  (h#h$e]r˂  (h	he]r̂  (hh�e]r͂  (h)heeej��  j��  ]r΂  (j�^  ]rς  (j�^  ]rЂ  (j�^  ]rт  (h	h�e]r҂  (hh�e]rӂ  (hhe]rԂ  (j�^  ]rՂ  (h	he]rւ  (hh�e]rׂ  (hhe]r؂  (j}w  ]rق  (h	h�e]rڂ  (hh�eeee]rۂ  (hhee]r܂  (h!]r݂  (h#h$e]rނ  (h	he]r߂  (hh�e]r��  (h)heeej΂  j΂  j΂  j΂  j΂  j΂  j΂  j΂  j΂  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r��  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r �  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej�  ]r�  (j�^  ]r�  (j�^  ]r	�  (j�^  ]r
�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r �  (j�^  ]r!�  (h	h�e]r"�  (hh�e]r#�  (hhe]r$�  (j}w  ]r%�  (h	h�e]r&�  (hh�eeee]r'�  (hhee]r(�  (h!]r)�  (h#h$e]r*�  (h	he]r+�  (hh�e]r,�  (h)heeej�  j�  j�  j�  ]r-�  (j�^  ]r.�  (j�^  ]r/�  (j�^  ]r0�  (h	h�e]r1�  (hh�e]r2�  (hhe]r3�  (j�^  ]r4�  (h	h�e]r5�  (hh�e]r6�  (hhe]r7�  (j}w  ]r8�  (h	h�e]r9�  (hh�eeee]r:�  (hhee]r;�  (h!]r<�  (h#h$e]r=�  (h	he]r>�  (hh�e]r?�  (h)heee]r@�  (j�^  ]rA�  (j�^  ]rB�  (j�^  ]rC�  (h	h�e]rD�  (hh�e]rE�  (hhe]rF�  (j�^  ]rG�  (h	h�e]rH�  (hh�e]rI�  (hhe]rJ�  (j}w  ]rK�  (h	h�e]rL�  (hh�eeee]rM�  (hhee]rN�  (h!]rO�  (h#h$e]rP�  (h	he]rQ�  (hh�e]rR�  (h)heeej@�  j@�  j@�  j@�  j@�  j@�  j@�  j@�  ]rS�  (j�^  ]rT�  (j�^  ]rU�  (j�^  ]rV�  (h	h�e]rW�  (hh�e]rX�  (hhe]rY�  (j�^  ]rZ�  (h	h�e]r[�  (hh�e]r\�  (hhe]r]�  (j}w  ]r^�  (h	h�e]r_�  (hh�eeee]r`�  (hhee]ra�  (h!]rb�  (h#h$e]rc�  (h	he]rd�  (hh�e]re�  (h)heeejS�  jS�  jS�  jS�  jS�  jS�  jS�  jS�  jS�  jS�  ]rf�  (j�^  ]rg�  (j�^  ]rh�  (j�^  ]ri�  (h	h�e]rj�  (hh�e]rk�  (hhe]rl�  (j�^  ]rm�  (h	h�e]rn�  (hh�e]ro�  (hhe]rp�  (j}w  ]rq�  (h	h�e]rr�  (hh�eeee]rs�  (hhee]rt�  (h!]ru�  (h#h$e]rv�  (h	he]rw�  (hh�e]rx�  (h)heee]ry�  (j�^  ]rz�  (j�^  ]r{�  (j�^  ]r|�  (h	h�e]r}�  (hh�e]r~�  (hhe]r�  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeejy�  jy�  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heee]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r  (h	he]rÃ  (hh�e]ră  (h)heeej��  j��  j��  j��  ]rŃ  (j�^  ]rƃ  (j�^  ]rǃ  (j�^  ]rȃ  (h	h�e]rɃ  (hh�e]rʃ  (hhe]r˃  (j�^  ]r̃  (h	he]r̓  (hh�e]r΃  (hhe]rσ  (j}w  ]rЃ  (h	h�e]rу  (hh�eeee]r҃  (hhee]rӃ  (h!]rԃ  (h#h$e]rՃ  (h	he]rփ  (hh�e]r׃  (h)heeejŃ  jŃ  ]r؃  (j�^  ]rك  (j�^  ]rڃ  (j�^  ]rۃ  (h	h�e]r܃  (hh�e]r݃  (hhe]rރ  (j�^  ]r߃  (h	he]r��  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r��  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej�  j�  j�  j�  j�  ]r��  (j�^  ]r��  (j�^  ]r �  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r	�  (h	h�e]r
�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej��  j��  j��  j��  j��  j��  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r �  (h#h$e]r!�  (h	he]r"�  (hh�e]r#�  (h)heeej�  j�  j�  ]r$�  (j�^  ]r%�  (j�^  ]r&�  (j�^  ]r'�  (h	h�e]r(�  (hh�e]r)�  (hhe]r*�  (j�^  ]r+�  (h	he]r,�  (hh�e]r-�  (hhe]r.�  (j}w  ]r/�  (h	h�e]r0�  (hh�eeee]r1�  (hhee]r2�  (h!]r3�  (h#h$e]r4�  (h	he]r5�  (hh�e]r6�  (h)heeej$�  j$�  j$�  ]r7�  (j�^  ]r8�  (j�^  ]r9�  (j�^  ]r:�  (h	h�e]r;�  (hh�e]r<�  (hhe]r=�  (j�^  ]r>�  (h	he]r?�  (hh�e]r@�  (hhe]rA�  (j}w  ]rB�  (h	h�e]rC�  (hh�eeee]rD�  (hhee]rE�  (h!]rF�  (h#h$e]rG�  (h	he]rH�  (hh�e]rI�  (h)heee]rJ�  (j�^  ]rK�  (j�^  ]rL�  (j�^  ]rM�  (h	h�e]rN�  (hh�e]rO�  (hhe]rP�  (j�^  ]rQ�  (h	he]rR�  (hh�e]rS�  (hhe]rT�  (j}w  ]rU�  (h	h�e]rV�  (hh�eeee]rW�  (hhee]rX�  (h!]rY�  (h#h$e]rZ�  (h	he]r[�  (hh�e]r\�  (h)heeejJ�  jJ�  ]r]�  (j�^  ]r^�  (j�^  ]r_�  (j�^  ]r`�  (h	h�e]ra�  (hh�e]rb�  (hhe]rc�  (j�^  ]rd�  (h	he]re�  (hh�e]rf�  (hhe]rg�  (j}w  ]rh�  (h	h�e]ri�  (hh�eeee]rj�  (hhee]rk�  (h!]rl�  (h#h$e]rm�  (h	he]rn�  (hh�e]ro�  (h)heeej]�  j]�  j]�  ]rp�  (j�^  ]rq�  (j�^  ]rr�  (j�^  ]rs�  (h	h�e]rt�  (hh�e]ru�  (hhe]rv�  (j�^  ]rw�  (h	he]rx�  (hh�e]ry�  (hhe]rz�  (j}w  ]r{�  (h	h�e]r|�  (hh�eeee]r}�  (hhee]r~�  (h!]r�  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeejp�  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r  (j�^  ]rÄ  (h	he]rĄ  (hh�e]rń  (hhe]rƄ  (j}w  ]rǄ  (h	h�e]rȄ  (hh�eeee]rɄ  (hhee]rʄ  (h!]r˄  (h#h$e]r̄  (h	he]r̈́  (hh�e]r΄  (h)heeej��  j��  j��  j��  j��  j��  ]rτ  (j�^  ]rЄ  (j�^  ]rф  (j�^  ]r҄  (h	h�e]rӄ  (hh�e]rԄ  (hhe]rՄ  (j�^  ]rք  (h	he]rׄ  (hh�e]r؄  (hhe]rل  (j}w  ]rڄ  (h	h�e]rۄ  (hh�eeee]r܄  (hhee]r݄  (h!]rބ  (h#h$e]r߄  (h	he]r��  (hh�e]r�  (h)heeejτ  jτ  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r��  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r �  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  ]r�  (j�^  ]r	�  (j�^  ]r
�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r �  (hhe]r!�  (j�^  ]r"�  (h	he]r#�  (hh�e]r$�  (hhe]r%�  (j}w  ]r&�  (h	h�e]r'�  (hh�eeee]r(�  (hhee]r)�  (h!]r*�  (h#h$e]r+�  (h	he]r,�  (hh�e]r-�  (h)heeej�  j�  j�  ]r.�  (j�^  ]r/�  (j�^  ]r0�  (j�^  ]r1�  (h	h�e]r2�  (hh�e]r3�  (hhe]r4�  (j�^  ]r5�  (h	he]r6�  (hh�e]r7�  (hhe]r8�  (j}w  ]r9�  (h	h�e]r:�  (hh�eeee]r;�  (hhee]r<�  (h!]r=�  (h#h$e]r>�  (h	he]r?�  (hh�e]r@�  (h)heeej.�  j.�  ]rA�  (j�^  ]rB�  (j�^  ]rC�  (j�^  ]rD�  (h	h�e]rE�  (hh�e]rF�  (hhe]rG�  (j�^  ]rH�  (h	he]rI�  (hh�e]rJ�  (hhe]rK�  (j}w  ]rL�  (h	h�e]rM�  (hh�eeee]rN�  (hhee]rO�  (h!]rP�  (h#h$e]rQ�  (h	he]rR�  (hh�e]rS�  (h)heeejA�  jA�  ]rT�  (j�^  ]rU�  (j�^  ]rV�  (j�^  ]rW�  (h	h�e]rX�  (hh�e]rY�  (hhe]rZ�  (j�^  ]r[�  (h	he]r\�  (hh�e]r]�  (hhe]r^�  (j}w  ]r_�  (h	h�e]r`�  (hh�eeee]ra�  (hhee]rb�  (h!]rc�  (h#h$e]rd�  (h	he]re�  (hh�e]rf�  (h)heeejT�  jT�  ]rg�  (j�^  ]rh�  (j�^  ]ri�  (j�^  ]rj�  (h	h�e]rk�  (hh�e]rl�  (hhe]rm�  (j�^  ]rn�  (h	he]ro�  (hh�e]rp�  (hhe]rq�  (j}w  ]rr�  (h	h�e]rs�  (hh�eeee]rt�  (hhee]ru�  (h!]rv�  (h#h$e]rw�  (h	he]rx�  (hh�e]ry�  (h)heee]rz�  (j�^  ]r{�  (j�^  ]r|�  (j�^  ]r}�  (h	h�e]r~�  (hh�e]r�  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeejz�  jz�  jz�  jz�  jz�  jz�  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r  (h#h$e]rÅ  (h	he]rą  (hh�e]rŅ  (h)heeej��  j��  ]rƅ  (j�^  ]rǅ  (j�^  ]rȅ  (j�^  ]rɅ  (h	h�e]rʅ  (hh�e]r˅  (hhe]r̅  (j�^  ]rͅ  (h	h�e]r΅  (hh�e]rυ  (hhe]rЅ  (j}w  ]rх  (h	h�e]r҅  (hh�eeee]rӅ  (hhee]rԅ  (h!]rՅ  (h#h$e]rօ  (h	he]rׅ  (hh�e]r؅  (h)heeejƅ  ]rم  (j�^  ]rڅ  (j�^  ]rۅ  (j�^  ]r܅  (h	h�e]r݅  (hh�e]rޅ  (hhe]r߅  (j�^  ]r��  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r��  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heee]r��  (j�^  ]r �  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r	�  (j}w  ]r
�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej��  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r �  (h!]r!�  (h#h$e]r"�  (h	he]r#�  (hh�e]r$�  (h)heeej�  j�  ]r%�  (j�^  ]r&�  (j�^  ]r'�  (j�^  ]r(�  (h	h�e]r)�  (hh�e]r*�  (hhe]r+�  (j�^  ]r,�  (h	h�e]r-�  (hh�e]r.�  (hhe]r/�  (j}w  ]r0�  (h	h�e]r1�  (hh�eeee]r2�  (hhee]r3�  (h!]r4�  (h#h$e]r5�  (h	he]r6�  (hh�e]r7�  (h)heeej%�  ]r8�  (j�^  ]r9�  (j�^  ]r:�  (j�^  ]r;�  (h	h�e]r<�  (hh�e]r=�  (hhe]r>�  (j�^  ]r?�  (h	h�e]r@�  (hh�e]rA�  (hhe]rB�  (j}w  ]rC�  (h	h�e]rD�  (hh�eeee]rE�  (hhee]rF�  (h!]rG�  (h#h$e]rH�  (h	he]rI�  (hh�e]rJ�  (h)heeej8�  ]rK�  (j�^  ]rL�  (j�^  ]rM�  (j�^  ]rN�  (h	h�e]rO�  (hh�e]rP�  (hhe]rQ�  (j�^  ]rR�  (h	h�e]rS�  (hh�e]rT�  (hhe]rU�  (j}w  ]rV�  (h	h�e]rW�  (hh�eeee]rX�  (hhee]rY�  (h!]rZ�  (h#h$e]r[�  (h	he]r\�  (hh�e]r]�  (h)heeejK�  jK�  jK�  jK�  ]r^�  (j�^  ]r_�  (j�^  ]r`�  (j�^  ]ra�  (h	h�e]rb�  (hh�e]rc�  (hhe]rd�  (j�^  ]re�  (h	h�e]rf�  (hh�e]rg�  (hhe]rh�  (j}w  ]ri�  (h	h�e]rj�  (hh�eeee]rk�  (hhee]rl�  (h!]rm�  (h#h$e]rn�  (h	he]ro�  (hh�e]rp�  (h)heeej^�  ]rq�  (j�^  ]rr�  (j�^  ]rs�  (j�^  ]rt�  (h	h�e]ru�  (hh�e]rv�  (hhe]rw�  (j�^  ]rx�  (h	h�e]ry�  (hh�e]rz�  (hhe]r{�  (j}w  ]r|�  (h	h�e]r}�  (hh�eeee]r~�  (hhee]r�  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeejq�  jq�  jq�  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heee]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r  (hhe]rÆ  (j�^  ]rĆ  (h	he]rņ  (hh�e]rƆ  (hhe]rǆ  (j}w  ]rȆ  (h	h�e]rɆ  (hh�eeee]rʆ  (hhee]rˆ  (h!]r̆  (h#h$e]r͆  (h	he]rΆ  (hh�e]rφ  (h)heeej��  j��  j��  j��  ]rІ  (j�^  ]rц  (j�^  ]r҆  (j�^  ]rӆ  (h	h�e]rԆ  (hh�e]rՆ  (hhe]rֆ  (j�^  ]r׆  (h	he]r؆  (hh�e]rن  (hhe]rچ  (j}w  ]rۆ  (h	h�e]r܆  (hh�eeee]r݆  (hhee]rކ  (h!]r߆  (h#h$e]r��  (h	he]r�  (hh�e]r�  (h)heeejІ  jІ  jІ  jІ  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r��  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r��  (h)heeej�  j�  j�  j�  j�  ]r��  (j�^  ]r��  (j�^  ]r��  (j�^  ]r��  (h	h�e]r��  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r �  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej��  ]r	�  (j�^  ]r
�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r�  (hh�e]r�  (hhe]r�  (j�^  ]r�  (h	he]r�  (hh�e]r�  (hhe]r�  (j}w  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej	�  j	�  j	�  j	�  j	�  j	�  j	�  j	�  j	�  ]r�  (j�^  ]r�  (j�^  ]r�  (j�^  ]r�  (h	h�e]r �  (hh�e]r!�  (hhe]r"�  (j�^  ]r#�  (h	he]r$�  (hh�e]r%�  (hhe]r&�  (j}w  ]r'�  (h	h�e]r(�  (hh�eeee]r)�  (hhee]r*�  (h!]r+�  (h#h$e]r,�  (h	he]r-�  (hh�e]r.�  (h)heeej�  j�  j�  j�  j�  j�  j�  ]r/�  (j�^  ]r0�  (j�^  ]r1�  (j�^  ]r2�  (h	h�e]r3�  (hh�e]r4�  (hhe]r5�  (j�^  ]r6�  (h	he]r7�  (hh�e]r8�  (hhe]r9�  (j}w  ]r:�  (h	h�e]r;�  (hh�eeee]r<�  (hhee]r=�  (h!]r>�  (h#h$e]r?�  (h	he]r@�  (hh�e]rA�  (h)heeej/�  ]rB�  (j�^  ]rC�  (j�^  ]rD�  (j�^  ]rE�  (h	h�e]rF�  (hh�e]rG�  (hhe]rH�  (j�^  ]rI�  (h	he]rJ�  (hh�e]rK�  (hhe]rL�  (j}w  ]rM�  (h	h�e]rN�  (hh�eeee]rO�  (hhee]rP�  (h!]rQ�  (h#h$e]rR�  (h	he]rS�  (hh�e]rT�  (h)heeejB�  jB�  ]rU�  (j�^  ]rV�  (j�^  ]rW�  (j�^  ]rX�  (h	h�e]rY�  (hh�e]rZ�  (hhe]r[�  (j�^  ]r\�  (h	he]r]�  (hh�e]r^�  (hhe]r_�  (j}w  ]r`�  (h	h�e]ra�  (hh�eeee]rb�  (hhee]rc�  (h!]rd�  (h#h$e]re�  (h	he]rf�  (hh�e]rg�  (h)heee]rh�  (j�^  ]ri�  (j�^  ]rj�  (j�^  ]rk�  (h	h�e]rl�  (hh�e]rm�  (hhe]rn�  (j�^  ]ro�  (h	he]rp�  (hh�e]rq�  (hhe]rr�  (j}w  ]rs�  (h	h�e]rt�  (hh�eeee]ru�  (hhee]rv�  (h!]rw�  (h#h$e]rx�  (h	he]ry�  (hh�e]rz�  (h)heee]r{�  (j�^  ]r|�  (j�^  ]r}�  (j�^  ]r~�  (h	h�e]r�  (hh�e]r��  (hhe]r��  (j�^  ]r��  (h	he]r��  (hh�e]r��  (hhe]r��  (j}w  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeee(j{�  e]r��  (]r��  (X   Normsr��  ]r��  (X   Oblr��  ]r��  (X   Movedr��  ]r��  (h	h
e]r��  (hX   anyr��  e]r��  (hhe]r��  (X   Movedr��  ]r��  (h	h
e]r��  (hX   circler��  e]r��  (hhe]r��  (X	   Next-Mover��  ]r��  (h	he]r��  (hX   triangler��  eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	X   anyr��  e]r��  (hX   triangler��  e]r��  (h)heeej��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hj��  e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hj��  e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hj��  eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j��  e]r��  (hh<e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r  (h	h
e]rÇ  (hj��  e]rć  (hhe]rŇ  (j��  ]rƇ  (h	h
e]rǇ  (hj��  e]rȇ  (hhe]rɇ  (j��  ]rʇ  (h	he]rˇ  (hj��  eeee]ṙ  (hhee]r͇  (h!]r·  (h#h$e]rχ  (h	h�e]rЇ  (hh<e]rч  (h)heeej��  ]r҇  (j��  ]rӇ  (j��  ]rԇ  (j��  ]rՇ  (h	h
e]rև  (hh�e]rׇ  (hhe]r؇  (j��  ]rه  (h	h
e]rڇ  (hj��  e]rۇ  (hhe]r܇  (j��  ]r݇  (h	he]rއ  (hj��  eeee]r߇  (hhee]r��  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)heeej҇  j҇  j҇  j҇  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hj��  e]r�  (hhe]r�  (j��  ]r��  (h	he]r�  (hj��  eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r��  (h	he]r��  (hh<e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r �  (hj��  e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hj��  eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r	�  (hh<e]r
�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hj��  e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hj��  eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r �  (j��  ]r!�  (h	h
e]r"�  (hh�e]r#�  (hhe]r$�  (j��  ]r%�  (h	h
e]r&�  (hj��  e]r'�  (hhe]r(�  (j��  ]r)�  (h	he]r*�  (hj��  eeee]r+�  (hhee]r,�  (h!]r-�  (h#h$e]r.�  (h	he]r/�  (hh�e]r0�  (h)heee]r1�  (j��  ]r2�  (j��  ]r3�  (j��  ]r4�  (h	h
e]r5�  (hh�e]r6�  (hhe]r7�  (j��  ]r8�  (h	h�e]r9�  (hj��  e]r:�  (hhe]r;�  (j��  ]r<�  (h	he]r=�  (hj��  eeee]r>�  (hhee]r?�  (h!]r@�  (h#h$e]rA�  (h	he]rB�  (hh�e]rC�  (h)heee]rD�  (j��  ]rE�  (j��  ]rF�  (j��  ]rG�  (h	h
e]rH�  (hh�e]rI�  (hhe]rJ�  (j��  ]rK�  (h	h�e]rL�  (hj��  e]rM�  (hhe]rN�  (j��  ]rO�  (h	he]rP�  (hj��  eeee]rQ�  (hhee]rR�  (h!]rS�  (h#h$e]rT�  (h	he]rU�  (hh�e]rV�  (h)heee]rW�  (j��  ]rX�  (j��  ]rY�  (j��  ]rZ�  (h	h
e]r[�  (hh�e]r\�  (hhe]r]�  (j��  ]r^�  (h	h�e]r_�  (hj��  e]r`�  (hhe]ra�  (j��  ]rb�  (h	he]rc�  (hj��  eeee]rd�  (hhee]re�  (h!]rf�  (h#h$e]rg�  (h	he]rh�  (hh�e]ri�  (h)heeejW�  ]rj�  (j��  ]rk�  (j��  ]rl�  (j��  ]rm�  (h	h
e]rn�  (hh�e]ro�  (hhe]rp�  (j��  ]rq�  (h	h�e]rr�  (hj��  e]rs�  (hhe]rt�  (j��  ]ru�  (h	he]rv�  (hj��  eeee]rw�  (hhee]rx�  (h!]ry�  (h#h$e]rz�  (h	h�e]r{�  (hh�e]r|�  (h)heee]r}�  (j��  ]r~�  (j��  ]r�  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r  (hj��  eeee]rÈ  (hhee]rĈ  (h!]rň  (h#h$e]rƈ  (h	h�e]rǈ  (hh�e]rȈ  (h)heee]rɈ  (j��  ]rʈ  (j��  ]rˈ  (j��  ]r̈  (h	h
e]r͈  (hh�e]rΈ  (hhe]rψ  (j��  ]rЈ  (h	h�e]rш  (hj��  e]r҈  (hhe]rӈ  (j��  ]rԈ  (h	h�e]rՈ  (hj��  eeee]rֈ  (hhee]r׈  (h!]r؈  (h#h$e]rو  (h	h�e]rڈ  (hh�e]rۈ  (h)heee]r܈  (j��  ]r݈  (j��  ]rވ  (j��  ]r߈  (h	h
e]r��  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hj��  e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hj��  eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r��  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r �  (hh<e]r�  (h)heeej�  j�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r	�  (h	h�e]r
�  (hj��  e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hj��  eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hj��  e]r�  (hhe]r�  (j��  ]r �  (h	h�e]r!�  (hj��  eeee]r"�  (hhee]r#�  (h!]r$�  (h#h$e]r%�  (h	j�  e]r&�  (hh<e]r'�  (h)heee]r(�  (j��  ]r)�  (j��  ]r*�  (j��  ]r+�  (h	h
e]r,�  (hh�e]r-�  (hhe]r.�  (j��  ]r/�  (h	h�e]r0�  (hj��  e]r1�  (hhe]r2�  (j��  ]r3�  (h	h�e]r4�  (hj��  eeee]r5�  (hhee]r6�  (h!]r7�  (h#h$e]r8�  (h	h
e]r9�  (hh<e]r:�  (h)heeej(�  j(�  j(�  j(�  j(�  j(�  ]r;�  (j��  ]r<�  (j��  ]r=�  (j��  ]r>�  (h	h
e]r?�  (hh�e]r@�  (hhe]rA�  (j��  ]rB�  (h	h�e]rC�  (hj��  e]rD�  (hhe]rE�  (j��  ]rF�  (h	h�e]rG�  (hj��  eeee]rH�  (hhee]rI�  (h!]rJ�  (h#h$e]rK�  (h	j�  e]rL�  (hh<e]rM�  (h)heeej;�  j;�  j;�  ]rN�  (j��  ]rO�  (j��  ]rP�  (j��  ]rQ�  (h	h
e]rR�  (hh�e]rS�  (hhe]rT�  (j��  ]rU�  (h	h�e]rV�  (hj��  e]rW�  (hhe]rX�  (j��  ]rY�  (h	h�e]rZ�  (hj��  eeee]r[�  (hhee]r\�  (h!]r]�  (h#h$e]r^�  (h	j�  e]r_�  (hh<e]r`�  (h)heeejN�  jN�  ]ra�  (j��  ]rb�  (j��  ]rc�  (j��  ]rd�  (h	h
e]re�  (hh�e]rf�  (hhe]rg�  (j��  ]rh�  (h	h�e]ri�  (hj��  e]rj�  (hhe]rk�  (j��  ]rl�  (h	h�e]rm�  (hj��  eeee]rn�  (hhee]ro�  (h!]rp�  (h#h$e]rq�  (h	j�  e]rr�  (hh<e]rs�  (h)heeeja�  ja�  ja�  ja�  ja�  ]rt�  (j��  ]ru�  (j��  ]rv�  (j��  ]rw�  (h	h
e]rx�  (hh�e]ry�  (hhe]rz�  (j��  ]r{�  (h	h�e]r|�  (hj��  e]r}�  (hhe]r~�  (j��  ]r�  (h	h�e]r��  (hj��  eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heeejt�  jt�  jt�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hj��  eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r  (j��  ]rÉ  (h	h
e]rĉ  (hh�e]rŉ  (hhe]rƉ  (j��  ]rǉ  (h	h�e]rȉ  (hj��  e]rɉ  (hhe]rʉ  (j��  ]rˉ  (h	he]r̉  (hj��  eeee]r͉  (hhee]rΉ  (h!]rω  (h#h$e]rЉ  (h	h�e]rщ  (hh�e]r҉  (h)heee]rӉ  (j��  ]rԉ  (j��  ]rՉ  (j��  ]r։  (h	h
e]r׉  (hh�e]r؉  (hhe]rى  (j��  ]rډ  (h	h�e]rۉ  (hj��  e]r܉  (hhe]r݉  (j��  ]rމ  (h	he]r߉  (hj��  eeee]r��  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hj��  e]r�  (hhe]r��  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r �  (h	h�e]r�  (hj��  e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r	�  (h	h�e]r
�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hj��  e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (j��  ]r �  (j��  ]r!�  (j��  ]r"�  (h	h
e]r#�  (hh�e]r$�  (hhe]r%�  (j��  ]r&�  (h	h�e]r'�  (hj��  e]r(�  (hhe]r)�  (j��  ]r*�  (h	he]r+�  (hh�eeee]r,�  (hhee]r-�  (h!]r.�  (h#h$e]r/�  (h	h�e]r0�  (hh�e]r1�  (h)heee]r2�  (j��  ]r3�  (j��  ]r4�  (j��  ]r5�  (h	h
e]r6�  (hh�e]r7�  (hhe]r8�  (j��  ]r9�  (h	h�e]r:�  (hj��  e]r;�  (hhe]r<�  (j��  ]r=�  (h	he]r>�  (hh�eeee]r?�  (hhee]r@�  (h!]rA�  (h#h$e]rB�  (h	h�e]rC�  (hh�e]rD�  (h)heee]rE�  (j��  ]rF�  (j��  ]rG�  (j��  ]rH�  (h	h
e]rI�  (hh�e]rJ�  (hhe]rK�  (j��  ]rL�  (h	h�e]rM�  (hj��  e]rN�  (hhe]rO�  (j��  ]rP�  (h	he]rQ�  (hh�eeee]rR�  (hhee]rS�  (h!]rT�  (h#h$e]rU�  (h	h�e]rV�  (hh�e]rW�  (h)heee]rX�  (j��  ]rY�  (j��  ]rZ�  (j��  ]r[�  (h	h
e]r\�  (hh<e]r]�  (hhe]r^�  (j��  ]r_�  (h	h�e]r`�  (hj��  e]ra�  (hhe]rb�  (j��  ]rc�  (h	he]rd�  (hh�eeee]re�  (hhee]rf�  (h!]rg�  (h#h$e]rh�  (h	h�e]ri�  (hh�e]rj�  (h)heeejX�  ]rk�  (j��  ]rl�  (j��  ]rm�  (j��  ]rn�  (h	h
e]ro�  (hh<e]rp�  (hhe]rq�  (j��  ]rr�  (h	h
e]rs�  (hj��  e]rt�  (hhe]ru�  (j��  ]rv�  (h	he]rw�  (hh�eeee]rx�  (hhee]ry�  (h!]rz�  (h#h$e]r{�  (h	h�e]r|�  (hh�e]r}�  (h)heeejk�  ]r~�  (j��  ]r�  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hj��  e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej~�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r  (h	he]rÊ  (hh�eeee]rĊ  (hhee]rŊ  (h!]rƊ  (h#h$e]rǊ  (h	h�e]rȊ  (hh�e]rɊ  (h)heeej��  j��  ]rʊ  (j��  ]rˊ  (j��  ]r̊  (j��  ]r͊  (h	h
e]rΊ  (hh<e]rϊ  (hhe]rЊ  (j��  ]rъ  (h	h
e]rҊ  (hh�e]rӊ  (hhe]rԊ  (j��  ]rՊ  (h	he]r֊  (hh�eeee]r׊  (hhee]r؊  (h!]rي  (h#h$e]rڊ  (h	h�e]rۊ  (hh�e]r܊  (h)heeejʊ  jʊ  ]r݊  (j��  ]rފ  (j��  ]rߊ  (j��  ]r��  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r��  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r �  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r	�  (j��  ]r
�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r �  (j��  ]r!�  (h	h�e]r"�  (hh�eeee]r#�  (hhee]r$�  (h!]r%�  (h#h$e]r&�  (h	h�e]r'�  (hh�e]r(�  (h)heee]r)�  (j��  ]r*�  (j��  ]r+�  (j��  ]r,�  (h	h�e]r-�  (hh<e]r.�  (hhe]r/�  (j��  ]r0�  (h	h
e]r1�  (hh�e]r2�  (hhe]r3�  (j��  ]r4�  (h	h�e]r5�  (hh�eeee]r6�  (hhee]r7�  (h!]r8�  (h#h$e]r9�  (h	h�e]r:�  (hh�e]r;�  (h)heeej)�  ]r<�  (j��  ]r=�  (j��  ]r>�  (j��  ]r?�  (h	h�e]r@�  (hh<e]rA�  (hhe]rB�  (j��  ]rC�  (h	h
e]rD�  (hh�e]rE�  (hhe]rF�  (j��  ]rG�  (h	h�e]rH�  (hh�eeee]rI�  (hhee]rJ�  (h!]rK�  (h#h$e]rL�  (h	h�e]rM�  (hh�e]rN�  (h)heee]rO�  (j��  ]rP�  (j��  ]rQ�  (j��  ]rR�  (h	h�e]rS�  (hh<e]rT�  (hhe]rU�  (j��  ]rV�  (h	h
e]rW�  (hh�e]rX�  (hhe]rY�  (j��  ]rZ�  (h	h�e]r[�  (hh�eeee]r\�  (hhee]r]�  (h!]r^�  (h#h$e]r_�  (h	h�e]r`�  (hh�e]ra�  (h)heee]rb�  (j��  ]rc�  (j��  ]rd�  (j��  ]re�  (h	h�e]rf�  (hh<e]rg�  (hhe]rh�  (j��  ]ri�  (h	h
e]rj�  (hh�e]rk�  (hhe]rl�  (j��  ]rm�  (h	h�e]rn�  (hh�eeee]ro�  (hhee]rp�  (h!]rq�  (h#h$e]rr�  (h	h�e]rs�  (hh�e]rt�  (h)heeejb�  jb�  ]ru�  (j��  ]rv�  (j��  ]rw�  (j��  ]rx�  (h	h�e]ry�  (hh<e]rz�  (hhe]r{�  (j��  ]r|�  (h	h
e]r}�  (hh�e]r~�  (hhe]r�  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeeju�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r  (j��  ]rË  (j��  ]rċ  (h	h�e]rŋ  (hh<e]rƋ  (hhe]rǋ  (j��  ]rȋ  (h	h
e]rɋ  (hh�e]rʋ  (hhe]rˋ  (j��  ]r̋  (h	he]r͋  (hh�eeee]r΋  (hhee]rϋ  (h!]rЋ  (h#h$e]rы  (h	h�e]rҋ  (hh�e]rӋ  (h)heeej��  j��  ]rԋ  (j��  ]rՋ  (j��  ]r֋  (j��  ]r׋  (h	h�e]r؋  (hh<e]rً  (hhe]rڋ  (j��  ]rۋ  (h	h
e]r܋  (hh�e]r݋  (hhe]rދ  (j��  ]rߋ  (h	he]r��  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r��  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r �  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r	�  (h#h$e]r
�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r �  (j��  ]r!�  (j��  ]r"�  (j��  ]r#�  (h	h�e]r$�  (hh<e]r%�  (hhe]r&�  (j��  ]r'�  (h	h
e]r(�  (hh�e]r)�  (hhe]r*�  (j��  ]r+�  (h	h�e]r,�  (hh�eeee]r-�  (hhee]r.�  (h!]r/�  (h#h$e]r0�  (h	h�e]r1�  (hh�e]r2�  (h)heeej �  ]r3�  (j��  ]r4�  (j��  ]r5�  (j��  ]r6�  (h	h�e]r7�  (hh<e]r8�  (hhe]r9�  (j��  ]r:�  (h	h
e]r;�  (hh�e]r<�  (hhe]r=�  (j��  ]r>�  (h	h�e]r?�  (hh�eeee]r@�  (hhee]rA�  (h!]rB�  (h#h$e]rC�  (h	h
e]rD�  (hh�e]rE�  (h)heeej3�  j3�  j3�  j3�  j3�  j3�  ]rF�  (j��  ]rG�  (j��  ]rH�  (j��  ]rI�  (h	h�e]rJ�  (hh<e]rK�  (hhe]rL�  (j��  ]rM�  (h	h
e]rN�  (hh�e]rO�  (hhe]rP�  (j��  ]rQ�  (h	h�e]rR�  (hh�eeee]rS�  (hhee]rT�  (h!]rU�  (h#h$e]rV�  (h	j�  e]rW�  (hh�e]rX�  (h)heeejF�  jF�  jF�  ]rY�  (j��  ]rZ�  (j��  ]r[�  (j��  ]r\�  (h	h�e]r]�  (hh<e]r^�  (hhe]r_�  (j��  ]r`�  (h	h
e]ra�  (hh�e]rb�  (hhe]rc�  (j��  ]rd�  (h	h�e]re�  (hh�eeee]rf�  (hhee]rg�  (h!]rh�  (h#h$e]ri�  (h	j�  e]rj�  (hh�e]rk�  (h)heee]rl�  (j��  ]rm�  (j��  ]rn�  (j��  ]ro�  (h	h�e]rp�  (hh<e]rq�  (hhe]rr�  (j��  ]rs�  (h	h
e]rt�  (hh�e]ru�  (hhe]rv�  (j��  ]rw�  (h	h�e]rx�  (hh�eeee]ry�  (hhee]rz�  (h!]r{�  (h#h$e]r|�  (h	j�  e]r}�  (hh<e]r~�  (h)heee]r�  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)heeej�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)h�eeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r  (j��  ]rÌ  (h	h�e]rČ  (hh�eeee]rŌ  (hhee]rƌ  (h!]rǌ  (h#h$e]rȌ  (h	j�  e]rɌ  (hh<e]rʌ  (h)h�eeej��  j��  j��  ]rˌ  (j��  ]ř  (j��  ]r͌  (j��  ]rΌ  (h	h�e]rό  (hh<e]rЌ  (hhe]rь  (j��  ]rҌ  (h	h
e]rӌ  (hh�e]rԌ  (hhe]rՌ  (j��  ]r֌  (h	h�e]r׌  (hh�eeee]r،  (hhee]rٌ  (h!]rڌ  (h#h$e]rی  (h	j�  e]r܌  (hh<e]r݌  (h)h�eee]rތ  (j��  ]rߌ  (j��  ]r��  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r��  (h)h�eeejތ  jތ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r �  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)h�eee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r	�  (hhe]r
�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)h�eeej�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r �  (hhe]r!�  (j��  ]r"�  (h	h�e]r#�  (hh�eeee]r$�  (hhee]r%�  (h!]r&�  (h#h$e]r'�  (h	j�  e]r(�  (hh<e]r)�  (h)h�eeej�  ]r*�  (j��  ]r+�  (j��  ]r,�  (j��  ]r-�  (h	h
e]r.�  (hh<e]r/�  (hhe]r0�  (j��  ]r1�  (h	h
e]r2�  (hh�e]r3�  (hhe]r4�  (j��  ]r5�  (h	h�e]r6�  (hh�eeee]r7�  (hhee]r8�  (h!]r9�  (h#h$e]r:�  (h	j�  e]r;�  (hh<e]r<�  (h)h�eee]r=�  (j��  ]r>�  (j��  ]r?�  (j��  ]r@�  (h	h
e]rA�  (hh<e]rB�  (hhe]rC�  (j��  ]rD�  (h	h
e]rE�  (hh�e]rF�  (hhe]rG�  (j��  ]rH�  (h	h�e]rI�  (hh�eeee]rJ�  (hhee]rK�  (h!]rL�  (h#h$e]rM�  (h	j�  e]rN�  (hh<e]rO�  (h)h�eee]rP�  (j��  ]rQ�  (j��  ]rR�  (j��  ]rS�  (h	h
e]rT�  (hh<e]rU�  (hhe]rV�  (j��  ]rW�  (h	h
e]rX�  (hh�e]rY�  (hhe]rZ�  (j��  ]r[�  (h	h�e]r\�  (hh�eeee]r]�  (hhee]r^�  (h!]r_�  (h#h$e]r`�  (h	j�  e]ra�  (hh�e]rb�  (h)h�eee]rc�  (j��  ]rd�  (j��  ]re�  (j��  ]rf�  (h	h�e]rg�  (hh<e]rh�  (hhe]ri�  (j��  ]rj�  (h	h
e]rk�  (hh�e]rl�  (hhe]rm�  (j��  ]rn�  (h	h�e]ro�  (hh�eeee]rp�  (hhee]rq�  (h!]rr�  (h#h$e]rs�  (h	j�  e]rt�  (hh�e]ru�  (h)h�eeejc�  jc�  jc�  jc�  jc�  jc�  ]rv�  (j��  ]rw�  (j��  ]rx�  (j��  ]ry�  (h	h�e]rz�  (hh<e]r{�  (hhe]r|�  (j��  ]r}�  (h	h
e]r~�  (hh�e]r�  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heeejv�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heee]r  (j��  ]rÍ  (j��  ]rč  (j��  ]rō  (h	h
e]rƍ  (hh<e]rǍ  (hhe]rȍ  (j��  ]rɍ  (h	h
e]rʍ  (hh�e]rˍ  (hhe]r̍  (j��  ]r͍  (h	h�e]r΍  (hh�eeee]rύ  (hhee]rЍ  (h!]rэ  (h#h$e]rҍ  (h	j�  e]rӍ  (hh�e]rԍ  (h)heeej  ]rՍ  (j��  ]r֍  (j��  ]r׍  (j��  ]r؍  (h	h
e]rٍ  (hh<e]rڍ  (hhe]rۍ  (j��  ]r܍  (h	h
e]rݍ  (hh�e]rލ  (hhe]rߍ  (j��  ]r��  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeejՍ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r��  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heeej�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r �  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r	�  (h!]r
�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r �  (h)heee]r!�  (j��  ]r"�  (j��  ]r#�  (j��  ]r$�  (h	h
e]r%�  (hh<e]r&�  (hhe]r'�  (j��  ]r(�  (h	h
e]r)�  (hh�e]r*�  (hhe]r+�  (j��  ]r,�  (h	h�e]r-�  (hh�eeee]r.�  (hhee]r/�  (h!]r0�  (h#h$e]r1�  (h	j�  e]r2�  (hh�e]r3�  (h)heee]r4�  (j��  ]r5�  (j��  ]r6�  (j��  ]r7�  (h	h
e]r8�  (hh<e]r9�  (hhe]r:�  (j��  ]r;�  (h	h
e]r<�  (hh�e]r=�  (hhe]r>�  (j��  ]r?�  (h	h�e]r@�  (hh�eeee]rA�  (hhee]rB�  (h!]rC�  (h#h$e]rD�  (h	he]rE�  (hh�e]rF�  (h)heee]rG�  (j��  ]rH�  (j��  ]rI�  (j��  ]rJ�  (h	h
e]rK�  (hh<e]rL�  (hhe]rM�  (j��  ]rN�  (h	h
e]rO�  (hh�e]rP�  (hhe]rQ�  (j��  ]rR�  (h	h�e]rS�  (hh�eeee]rT�  (hhee]rU�  (h!]rV�  (h#h$e]rW�  (h	he]rX�  (hh�e]rY�  (h)heeejG�  ]rZ�  (j��  ]r[�  (j��  ]r\�  (j��  ]r]�  (h	h
e]r^�  (hh<e]r_�  (hhe]r`�  (j��  ]ra�  (h	h
e]rb�  (hh�e]rc�  (hhe]rd�  (j��  ]re�  (h	h�e]rf�  (hh�eeee]rg�  (hhee]rh�  (h!]ri�  (h#h$e]rj�  (h	j�  e]rk�  (hh�e]rl�  (h)heee]rm�  (j��  ]rn�  (j��  ]ro�  (j��  ]rp�  (h	h
e]rq�  (hh<e]rr�  (hhe]rs�  (j��  ]rt�  (h	h
e]ru�  (hh�e]rv�  (hhe]rw�  (j��  ]rx�  (h	he]ry�  (hh�eeee]rz�  (hhee]r{�  (h!]r|�  (h#h$e]r}�  (h	j�  e]r~�  (hh�e]r�  (h)heeejm�  jm�  jm�  jm�  jm�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh<e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh<e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh<e]r��  (h)heeej��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r  (hhe]rÎ  (j��  ]rĎ  (h	he]rŎ  (hh�eeee]rƎ  (hhee]rǎ  (h!]rȎ  (h#h$e]rɎ  (h	he]rʎ  (hh<e]rˎ  (h)heee]r̎  (j��  ]r͎  (j��  ]rΎ  (j��  ]rώ  (h	h
e]rЎ  (hh<e]rю  (hhe]rҎ  (j��  ]rӎ  (h	h
e]rԎ  (hh�e]rՎ  (hhe]r֎  (j��  ]r׎  (h	he]r؎  (hh�eeee]rَ  (hhee]rڎ  (h!]rێ  (h#h$e]r܎  (h	he]rݎ  (hh<e]rގ  (h)heeej̎  j̎  j̎  j̎  ]rߎ  (j��  ]r��  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r��  (hh<e]r�  (h)heeejߎ  jߎ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r �  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r	�  (hh<e]r
�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r �  (hh�e]r!�  (hhe]r"�  (j��  ]r#�  (h	he]r$�  (hh�eeee]r%�  (hhee]r&�  (h!]r'�  (h#h$e]r(�  (h	he]r)�  (hh<e]r*�  (h)heee]r+�  (j��  ]r,�  (j��  ]r-�  (j��  ]r.�  (h	h
e]r/�  (hh<e]r0�  (hhe]r1�  (j��  ]r2�  (h	h
e]r3�  (hh�e]r4�  (hhe]r5�  (j��  ]r6�  (h	he]r7�  (hh�eeee]r8�  (hhee]r9�  (h!]r:�  (h#h$e]r;�  (h	he]r<�  (hh<e]r=�  (h)heee]r>�  (j��  ]r?�  (j��  ]r@�  (j��  ]rA�  (h	h
e]rB�  (hh<e]rC�  (hhe]rD�  (j��  ]rE�  (h	h
e]rF�  (hh�e]rG�  (hhe]rH�  (j��  ]rI�  (h	he]rJ�  (hh�eeee]rK�  (hhee]rL�  (h!]rM�  (h#h$e]rN�  (h	he]rO�  (hh<e]rP�  (h)heeej>�  ]rQ�  (j��  ]rR�  (j��  ]rS�  (j��  ]rT�  (h	h
e]rU�  (hh<e]rV�  (hhe]rW�  (j��  ]rX�  (h	h
e]rY�  (hh�e]rZ�  (hhe]r[�  (j��  ]r\�  (h	he]r]�  (hh�eeee]r^�  (hhee]r_�  (h!]r`�  (h#h$e]ra�  (h	h
e]rb�  (hh<e]rc�  (h)heee]rd�  (j��  ]re�  (j��  ]rf�  (j��  ]rg�  (h	h
e]rh�  (hh<e]ri�  (hhe]rj�  (j��  ]rk�  (h	h
e]rl�  (hh�e]rm�  (hhe]rn�  (j��  ]ro�  (h	he]rp�  (hh�eeee]rq�  (hhee]rr�  (h!]rs�  (h#h$e]rt�  (h	h
e]ru�  (hh<e]rv�  (h)heeejd�  jd�  ]rw�  (j��  ]rx�  (j��  ]ry�  (j��  ]rz�  (h	h
e]r{�  (hh<e]r|�  (hhe]r}�  (j��  ]r~�  (h	h
e]r�  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh<e]r��  (h)heeejw�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r  (h)heeej��  j��  ]rÏ  (j��  ]rď  (j��  ]rŏ  (j��  ]rƏ  (h	h
e]rǏ  (hh<e]rȏ  (hhe]rɏ  (j��  ]rʏ  (h	h
e]rˏ  (hh�e]ȑ  (hhe]r͏  (j��  ]rΏ  (h	he]rϏ  (hh�eeee]rЏ  (hhee]rя  (h!]rҏ  (h#h$e]rӏ  (h	h
e]rԏ  (hh�e]rՏ  (h)heeejÏ  ]r֏  (j��  ]r׏  (j��  ]r؏  (j��  ]rُ  (h	h
e]rڏ  (hh<e]rۏ  (hhe]r܏  (j��  ]rݏ  (h	h
e]rޏ  (hh�e]rߏ  (hhe]r��  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r��  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)h�eee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r �  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r	�  (hhee]r
�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eeej��  j��  j��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r �  (hh�e]r!�  (h)h�eeej�  j�  ]r"�  (j��  ]r#�  (j��  ]r$�  (j��  ]r%�  (h	h
e]r&�  (hh<e]r'�  (hhe]r(�  (j��  ]r)�  (h	h
e]r*�  (hh�e]r+�  (hhe]r,�  (j��  ]r-�  (h	he]r.�  (hh�eeee]r/�  (hhee]r0�  (h!]r1�  (h#h$e]r2�  (h	h
e]r3�  (hh�e]r4�  (h)h�eee]r5�  (j��  ]r6�  (j��  ]r7�  (j��  ]r8�  (h	h
e]r9�  (hh<e]r:�  (hhe]r;�  (j��  ]r<�  (h	h
e]r=�  (hh�e]r>�  (hhe]r?�  (j��  ]r@�  (h	he]rA�  (hh�eeee]rB�  (hhee]rC�  (h!]rD�  (h#h$e]rE�  (h	h
e]rF�  (hh�e]rG�  (h)h�eeej5�  j5�  ]rH�  (j��  ]rI�  (j��  ]rJ�  (j��  ]rK�  (h	h
e]rL�  (hh<e]rM�  (hhe]rN�  (j��  ]rO�  (h	h
e]rP�  (hh�e]rQ�  (hhe]rR�  (j��  ]rS�  (h	he]rT�  (hh�eeee]rU�  (hhee]rV�  (h!]rW�  (h#h$e]rX�  (h	h
e]rY�  (hh�e]rZ�  (h)heee]r[�  (j��  ]r\�  (j��  ]r]�  (j��  ]r^�  (h	h
e]r_�  (hh<e]r`�  (hhe]ra�  (j��  ]rb�  (h	h
e]rc�  (hh�e]rd�  (hhe]re�  (j��  ]rf�  (h	he]rg�  (hh�eeee]rh�  (hhee]ri�  (h!]rj�  (h#h$e]rk�  (h	h
e]rl�  (hh�e]rm�  (h)heee]rn�  (j��  ]ro�  (j��  ]rp�  (j��  ]rq�  (h	h
e]rr�  (hh<e]rs�  (hhe]rt�  (j��  ]ru�  (h	h
e]rv�  (hh�e]rw�  (hhe]rx�  (j��  ]ry�  (h	he]rz�  (hh�eeee]r{�  (hhee]r|�  (h!]r}�  (h#h$e]r~�  (h	h
e]r�  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)h�eeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r  (hh<e]rÐ  (hhe]rĐ  (j��  ]rŐ  (h	he]rƐ  (hh�eeee]rǐ  (hhee]rȐ  (h!]rɐ  (h#h$e]rʐ  (h	j�  e]rː  (hh�e]r̐  (h)heee]r͐  (j��  ]rΐ  (j��  ]rϐ  (j��  ]rА  (h	h
e]rѐ  (hh<e]rҐ  (hhe]rӐ  (j��  ]rԐ  (h	h
e]rՐ  (hh<e]r֐  (hhe]rא  (j��  ]rؐ  (h	he]rِ  (hh�eeee]rڐ  (hhee]rې  (h!]rܐ  (h#h$e]rݐ  (h	j�  e]rސ  (hh�e]rߐ  (h)heeej͐  j͐  j͐  ]r��  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej��  ]r�  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r �  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r	�  (h	h
e]r
�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r �  (h	h�e]r!�  (hh<e]r"�  (hhe]r#�  (j��  ]r$�  (h	he]r%�  (hh�eeee]r&�  (hhee]r'�  (h!]r(�  (h#h$e]r)�  (h	j�  e]r*�  (hh<e]r+�  (h)heeej�  ]r,�  (j��  ]r-�  (j��  ]r.�  (j��  ]r/�  (h	h
e]r0�  (hh<e]r1�  (hhe]r2�  (j��  ]r3�  (h	h�e]r4�  (hh<e]r5�  (hhe]r6�  (j��  ]r7�  (h	he]r8�  (hh�eeee]r9�  (hhee]r:�  (h!]r;�  (h#h$e]r<�  (h	h
e]r=�  (hh<e]r>�  (h)heee]r?�  (j��  ]r@�  (j��  ]rA�  (j��  ]rB�  (h	h
e]rC�  (hh<e]rD�  (hhe]rE�  (j��  ]rF�  (h	h�e]rG�  (hh<e]rH�  (hhe]rI�  (j��  ]rJ�  (h	he]rK�  (hh�eeee]rL�  (hhee]rM�  (h!]rN�  (h#h$e]rO�  (h	h
e]rP�  (hh<e]rQ�  (h)heee]rR�  (j��  ]rS�  (j��  ]rT�  (j��  ]rU�  (h	h
e]rV�  (hh<e]rW�  (hhe]rX�  (j��  ]rY�  (h	h�e]rZ�  (hh<e]r[�  (hhe]r\�  (j��  ]r]�  (h	he]r^�  (hh�eeee]r_�  (hhee]r`�  (h!]ra�  (h#h$e]rb�  (h	h
e]rc�  (hh<e]rd�  (h)heee]re�  (j��  ]rf�  (j��  ]rg�  (j��  ]rh�  (h	h
e]ri�  (hh<e]rj�  (hhe]rk�  (j��  ]rl�  (h	h�e]rm�  (hh<e]rn�  (hhe]ro�  (j��  ]rp�  (h	he]rq�  (hh�eeee]rr�  (hhee]rs�  (h!]rt�  (h#h$e]ru�  (h	h
e]rv�  (hh<e]rw�  (h)heeeje�  ]rx�  (j��  ]ry�  (j��  ]rz�  (j��  ]r{�  (h	h
e]r|�  (hh<e]r}�  (hhe]r~�  (j��  ]r�  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh<e]r��  (h)heeejx�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh<e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh<e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r  (hh�e]rÑ  (h)heeej��  j��  j��  ]rđ  (j��  ]rő  (j��  ]rƑ  (j��  ]rǑ  (h	h
e]rȑ  (hh<e]rɑ  (hhe]rʑ  (j��  ]rˑ  (h	h�e]ȓ  (hh<e]r͑  (hhe]rΑ  (j��  ]rϑ  (h	he]rБ  (hh�eeee]rё  (hhee]rґ  (h!]rӑ  (h#h$e]rԑ  (h	j�  e]rՑ  (hh�e]r֑  (h)h�eeejđ  ]rב  (j��  ]rؑ  (j��  ]rّ  (j��  ]rڑ  (h	h
e]rۑ  (hh<e]rܑ  (hhe]rݑ  (j��  ]rޑ  (h	h�e]rߑ  (hh<e]r��  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)h�eeejב  jב  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)h�eeej�  j�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r �  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	he]r	�  (hh�eeee]r
�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)h�eee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r �  (h	j�  e]r!�  (hh<e]r"�  (h)h�eee]r#�  (j��  ]r$�  (j��  ]r%�  (j��  ]r&�  (h	h
e]r'�  (hh<e]r(�  (hhe]r)�  (j��  ]r*�  (h	h�e]r+�  (hh<e]r,�  (hhe]r-�  (j��  ]r.�  (h	he]r/�  (hh�eeee]r0�  (hhee]r1�  (h!]r2�  (h#h$e]r3�  (h	j�  e]r4�  (hh<e]r5�  (h)h�eee]r6�  (j��  ]r7�  (j��  ]r8�  (j��  ]r9�  (h	h
e]r:�  (hh<e]r;�  (hhe]r<�  (j��  ]r=�  (h	h�e]r>�  (hh<e]r?�  (hhe]r@�  (j��  ]rA�  (h	he]rB�  (hh�eeee]rC�  (hhee]rD�  (h!]rE�  (h#h$e]rF�  (h	j�  e]rG�  (hh<e]rH�  (h)h�eeej6�  j6�  ]rI�  (j��  ]rJ�  (j��  ]rK�  (j��  ]rL�  (h	h
e]rM�  (hh<e]rN�  (hhe]rO�  (j��  ]rP�  (h	h�e]rQ�  (hh<e]rR�  (hhe]rS�  (j��  ]rT�  (h	he]rU�  (hh�eeee]rV�  (hhee]rW�  (h!]rX�  (h#h$e]rY�  (h	j�  e]rZ�  (hh<e]r[�  (h)h�eeejI�  jI�  ]r\�  (j��  ]r]�  (j��  ]r^�  (j��  ]r_�  (h	h
e]r`�  (hh<e]ra�  (hhe]rb�  (j��  ]rc�  (h	h�e]rd�  (hh<e]re�  (hhe]rf�  (j��  ]rg�  (h	he]rh�  (hh�eeee]ri�  (hhee]rj�  (h!]rk�  (h#h$e]rl�  (h	j�  e]rm�  (hh<e]rn�  (h)h�eee]ro�  (j��  ]rp�  (j��  ]rq�  (j��  ]rr�  (h	h
e]rs�  (hh<e]rt�  (hhe]ru�  (j��  ]rv�  (h	h�e]rw�  (hh<e]rx�  (hhe]ry�  (j��  ]rz�  (h	he]r{�  (hh�eeee]r|�  (hhee]r}�  (h!]r~�  (h#h$e]r�  (h	j�  e]r��  (hh<e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r  (h	h�e]rÒ  (hh<e]rĒ  (hhe]rŒ  (j��  ]rƒ  (h	he]rǒ  (hh�eeee]rȒ  (hhee]rɒ  (h!]rʒ  (h#h$e]r˒  (h	j�  e]r̒  (hh<e]r͒  (h)heee]rΒ  (j��  ]rϒ  (j��  ]rВ  (j��  ]rђ  (h	h
e]rҒ  (hh<e]rӒ  (hhe]rԒ  (j��  ]rՒ  (h	h�e]r֒  (hh<e]rג  (hhe]rؒ  (j��  ]rْ  (h	he]rڒ  (hh�eeee]rے  (hhee]rܒ  (h!]rݒ  (h#h$e]rޒ  (h	j�  e]rߒ  (hh<e]r��  (h)heeejΒ  jΒ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r �  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r	�  (j��  ]r
�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r �  (j��  ]r!�  (h	h�e]r"�  (hh<e]r#�  (hhe]r$�  (j��  ]r%�  (h	he]r&�  (hh�eeee]r'�  (hhee]r(�  (h!]r)�  (h#h$e]r*�  (h	j�  e]r+�  (hh�e]r,�  (h)heee]r-�  (j��  ]r.�  (j��  ]r/�  (j��  ]r0�  (h	h
e]r1�  (hh<e]r2�  (hhe]r3�  (j��  ]r4�  (h	h
e]r5�  (hh<e]r6�  (hhe]r7�  (j��  ]r8�  (h	he]r9�  (hh�eeee]r:�  (hhee]r;�  (h!]r<�  (h#h$e]r=�  (h	j�  e]r>�  (hh�e]r?�  (h)heeej-�  j-�  j-�  j-�  j-�  j-�  j-�  ]r@�  (j��  ]rA�  (j��  ]rB�  (j��  ]rC�  (h	h
e]rD�  (hh<e]rE�  (hhe]rF�  (j��  ]rG�  (h	h
e]rH�  (hh<e]rI�  (hhe]rJ�  (j��  ]rK�  (h	he]rL�  (hh�eeee]rM�  (hhee]rN�  (h!]rO�  (h#h$e]rP�  (h	j�  e]rQ�  (hh�e]rR�  (h)heeej@�  ]rS�  (j��  ]rT�  (j��  ]rU�  (j��  ]rV�  (h	h
e]rW�  (hh<e]rX�  (hhe]rY�  (j��  ]rZ�  (h	h
e]r[�  (hh<e]r\�  (hhe]r]�  (j��  ]r^�  (h	he]r_�  (hh�eeee]r`�  (hhee]ra�  (h!]rb�  (h#h$e]rc�  (h	j�  e]rd�  (hh�e]re�  (h)heee]rf�  (j��  ]rg�  (j��  ]rh�  (j��  ]ri�  (h	h
e]rj�  (hh<e]rk�  (hhe]rl�  (j��  ]rm�  (h	h
e]rn�  (hh<e]ro�  (hhe]rp�  (j��  ]rq�  (h	he]rr�  (hh�eeee]rs�  (hhee]rt�  (h!]ru�  (h#h$e]rv�  (h	j�  e]rw�  (hh�e]rx�  (h)heeejf�  ]ry�  (j��  ]rz�  (j��  ]r{�  (j��  ]r|�  (h	h
e]r}�  (hh<e]r~�  (hhe]r�  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r  (h	j�  e]rÓ  (hh�e]rē  (h)heeej��  j��  j��  ]rœ  (j��  ]rƓ  (j��  ]rǓ  (j��  ]rȓ  (h	h
e]rɓ  (hh<e]rʓ  (hhe]r˓  (j��  ]r̓  (h	h
e]r͓  (hh<e]rΓ  (hhe]rϓ  (j��  ]rГ  (h	h�e]rѓ  (hh�eeee]rғ  (hhee]rӓ  (h!]rԓ  (h#h$e]rՓ  (h	he]r֓  (hh�e]rד  (h)heee]rؓ  (j��  ]rٓ  (j��  ]rړ  (j��  ]rۓ  (h	h
e]rܓ  (hh<e]rݓ  (hhe]rޓ  (j��  ]rߓ  (h	h
e]r��  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeejؓ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r �  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r	�  (h	h�e]r
�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)h�eee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r �  (h#h$e]r!�  (h	he]r"�  (hh<e]r#�  (h)h�eeej�  ]r$�  (j��  ]r%�  (j��  ]r&�  (j��  ]r'�  (h	h
e]r(�  (hh<e]r)�  (hhe]r*�  (j��  ]r+�  (h	h
e]r,�  (hh<e]r-�  (hhe]r.�  (j��  ]r/�  (h	h�e]r0�  (hh�eeee]r1�  (hhee]r2�  (h!]r3�  (h#h$e]r4�  (h	he]r5�  (hh<e]r6�  (h)heeej$�  ]r7�  (j��  ]r8�  (j��  ]r9�  (j��  ]r:�  (h	h
e]r;�  (hh<e]r<�  (hhe]r=�  (j��  ]r>�  (h	h
e]r?�  (hh<e]r@�  (hhe]rA�  (j��  ]rB�  (h	h�e]rC�  (hh�eeee]rD�  (hhee]rE�  (h!]rF�  (h#h$e]rG�  (h	h�e]rH�  (hh�e]rI�  (h)heeej7�  ]rJ�  (j��  ]rK�  (j��  ]rL�  (j��  ]rM�  (h	h
e]rN�  (hh<e]rO�  (hhe]rP�  (j��  ]rQ�  (h	h
e]rR�  (hh<e]rS�  (hhe]rT�  (j��  ]rU�  (h	h�e]rV�  (hh�eeee]rW�  (hhee]rX�  (h!]rY�  (h#h$e]rZ�  (h	h�e]r[�  (hh�e]r\�  (h)heee]r]�  (j��  ]r^�  (j��  ]r_�  (j��  ]r`�  (h	h
e]ra�  (hh<e]rb�  (hhe]rc�  (j��  ]rd�  (h	h
e]re�  (hh<e]rf�  (hhe]rg�  (j��  ]rh�  (h	h�e]ri�  (hh�eeee]rj�  (hhee]rk�  (h!]rl�  (h#h$e]rm�  (h	h�e]rn�  (hh�e]ro�  (h)heeej]�  ]rp�  (j��  ]rq�  (j��  ]rr�  (j��  ]rs�  (h	h
e]rt�  (hh<e]ru�  (hhe]rv�  (j��  ]rw�  (h	h
e]rx�  (hh<e]ry�  (hhe]rz�  (j��  ]r{�  (h	h�e]r|�  (hh�eeee]r}�  (hhee]r~�  (h!]r�  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r  (j��  ]rÔ  (h	h
e]rĔ  (hh<e]rŔ  (hhe]rƔ  (j��  ]rǔ  (h	h�e]rȔ  (hh�eeee]rɔ  (hhee]rʔ  (h!]r˔  (h#h$e]r̔  (h	h
e]r͔  (hh�e]rΔ  (h)heeej��  j��  j��  ]rϔ  (j��  ]rД  (j��  ]rє  (j��  ]rҔ  (h	h
e]rӔ  (hh�e]rԔ  (hhe]rՔ  (j��  ]r֔  (h	h
e]rה  (hh<e]rؔ  (hhe]rٔ  (j��  ]rڔ  (h	h�e]r۔  (hh�eeee]rܔ  (hhee]rݔ  (h!]rޔ  (h#h$e]rߔ  (h	h
e]r��  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r �  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heeej��  ]r�  (j��  ]r	�  (j��  ]r
�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r �  (hhe]r!�  (j��  ]r"�  (h	h
e]r#�  (hh<e]r$�  (hhe]r%�  (j��  ]r&�  (h	h�e]r'�  (hh�eeee]r(�  (hhee]r)�  (h!]r*�  (h#h$e]r+�  (h	h
e]r,�  (hh�e]r-�  (h)heee]r.�  (j��  ]r/�  (j��  ]r0�  (j��  ]r1�  (h	h
e]r2�  (hh<e]r3�  (hhe]r4�  (j��  ]r5�  (h	h
e]r6�  (hh<e]r7�  (hhe]r8�  (j��  ]r9�  (h	h�e]r:�  (hh�eeee]r;�  (hhee]r<�  (h!]r=�  (h#h$e]r>�  (h	h
e]r?�  (hh�e]r@�  (h)heeej.�  j.�  j.�  j.�  j.�  j.�  ]rA�  (j��  ]rB�  (j��  ]rC�  (j��  ]rD�  (h	h
e]rE�  (hh<e]rF�  (hhe]rG�  (j��  ]rH�  (h	h
e]rI�  (hh�e]rJ�  (hhe]rK�  (j��  ]rL�  (h	h�e]rM�  (hh�eeee]rN�  (hhee]rO�  (h!]rP�  (h#h$e]rQ�  (h	h
e]rR�  (hh�e]rS�  (h)heeejA�  jA�  jA�  jA�  ]rT�  (j��  ]rU�  (j��  ]rV�  (j��  ]rW�  (h	h
e]rX�  (hh<e]rY�  (hhe]rZ�  (j��  ]r[�  (h	h
e]r\�  (hh�e]r]�  (hhe]r^�  (j��  ]r_�  (h	h�e]r`�  (hh�eeee]ra�  (hhee]rb�  (h!]rc�  (h#h$e]rd�  (h	h
e]re�  (hh�e]rf�  (h)heee]rg�  (j��  ]rh�  (j��  ]ri�  (j��  ]rj�  (h	h
e]rk�  (hh<e]rl�  (hhe]rm�  (j��  ]rn�  (h	h
e]ro�  (hh�e]rp�  (hhe]rq�  (j��  ]rr�  (h	h�e]rs�  (hh�eeee]rt�  (hhee]ru�  (h!]rv�  (h#h$e]rw�  (h	h
e]rx�  (hh�e]ry�  (h)heee]rz�  (j��  ]r{�  (j��  ]r|�  (j��  ]r}�  (h	h
e]r~�  (hh<e]r�  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r  (h#h$e]rÕ  (h	j�  e]rĕ  (hh�e]rŕ  (h)heeej��  j��  ]rƕ  (j��  ]rǕ  (j��  ]rȕ  (j��  ]rɕ  (h	h�e]rʕ  (hh<e]r˕  (hhe]r̕  (j��  ]r͕  (h	h
e]rΕ  (hh�e]rϕ  (hhe]rЕ  (j��  ]rѕ  (h	h�e]rҕ  (hh�eeee]rӕ  (hhee]rԕ  (h!]rՕ  (h#h$e]r֕  (h	j�  e]rו  (hh�e]rؕ  (h)heee]rٕ  (j��  ]rڕ  (j��  ]rە  (j��  ]rܕ  (h	h�e]rݕ  (hh<e]rޕ  (hhe]rߕ  (j��  ]r��  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r �  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r	�  (j��  ]r
�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r �  (h!]r!�  (h#h$e]r"�  (h	h�e]r#�  (hh�e]r$�  (h)heeej�  j�  j�  j�  ]r%�  (j��  ]r&�  (j��  ]r'�  (j��  ]r(�  (h	h�e]r)�  (hh<e]r*�  (hhe]r+�  (j��  ]r,�  (h	h
e]r-�  (hh�e]r.�  (hhe]r/�  (j��  ]r0�  (h	h�e]r1�  (hh�eeee]r2�  (hhee]r3�  (h!]r4�  (h#h$e]r5�  (h	h
e]r6�  (hh�e]r7�  (h)h�eeej%�  j%�  ]r8�  (j��  ]r9�  (j��  ]r:�  (j��  ]r;�  (h	h�e]r<�  (hh<e]r=�  (hhe]r>�  (j��  ]r?�  (h	h
e]r@�  (hh�e]rA�  (hhe]rB�  (j��  ]rC�  (h	h�e]rD�  (hh�eeee]rE�  (hhee]rF�  (h!]rG�  (h#h$e]rH�  (h	h
e]rI�  (hh�e]rJ�  (h)h�eee]rK�  (j��  ]rL�  (j��  ]rM�  (j��  ]rN�  (h	h�e]rO�  (hh<e]rP�  (hhe]rQ�  (j��  ]rR�  (h	h
e]rS�  (hh�e]rT�  (hhe]rU�  (j��  ]rV�  (h	h�e]rW�  (hh�eeee]rX�  (hhee]rY�  (h!]rZ�  (h#h$e]r[�  (h	j�  e]r\�  (hh�e]r]�  (h)h�eeejK�  ]r^�  (j��  ]r_�  (j��  ]r`�  (j��  ]ra�  (h	h�e]rb�  (hh<e]rc�  (hhe]rd�  (j��  ]re�  (h	h
e]rf�  (hh�e]rg�  (hhe]rh�  (j��  ]ri�  (h	h�e]rj�  (hh�eeee]rk�  (hhee]rl�  (h!]rm�  (h#h$e]rn�  (h	j�  e]ro�  (hh�e]rp�  (h)h�eeej^�  j^�  ]rq�  (j��  ]rr�  (j��  ]rs�  (j��  ]rt�  (h	h�e]ru�  (hh<e]rv�  (hhe]rw�  (j��  ]rx�  (h	h
e]ry�  (hh�e]rz�  (hhe]r{�  (j��  ]r|�  (h	h�e]r}�  (hh�eeee]r~�  (hhee]r�  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)h�eeejq�  jq�  jq�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)h�eeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (X	   Next-Mover��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)h�eee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)h�eee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r  (hh<e]rÖ  (hhe]rĖ  (j��  ]rŖ  (h	h
e]rƖ  (hh�e]rǖ  (hhe]rȖ  (j��  ]rɖ  (h	he]rʖ  (hh�eeee]r˖  (hhee]r̖  (h!]r͖  (h#h$e]rΖ  (h	h
e]rϖ  (hh�e]rЖ  (h)heeej��  j��  ]rі  (j��  ]rҖ  (j��  ]rӖ  (j��  ]rԖ  (h	h�e]rՖ  (hh<e]r֖  (hhe]rז  (j��  ]rؖ  (h	h
e]rٖ  (hh�e]rږ  (hhe]rۖ  (j��  ]rܖ  (h	he]rݖ  (hh�eeee]rޖ  (hhee]rߖ  (h!]r��  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeejі  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heeej�  j�  j�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r �  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r	�  (h)heeej��  j��  j��  ]r
�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh�e]r�  (h)heeej
�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r �  (h	h
e]r!�  (hh<e]r"�  (hhe]r#�  (j��  ]r$�  (h	h
e]r%�  (hh�e]r&�  (hhe]r'�  (j��  ]r(�  (h	he]r)�  (hh�eeee]r*�  (hhee]r+�  (h!]r,�  (h#h$e]r-�  (h	j�  e]r.�  (hh�e]r/�  (h)heee]r0�  (j��  ]r1�  (j��  ]r2�  (j��  ]r3�  (h	h
e]r4�  (hh<e]r5�  (hhe]r6�  (j��  ]r7�  (h	h
e]r8�  (hh�e]r9�  (hhe]r:�  (j��  ]r;�  (h	he]r<�  (hh�eeee]r=�  (hhee]r>�  (h!]r?�  (h#h$e]r@�  (h	j�  e]rA�  (hh�e]rB�  (h)heeej0�  ]rC�  (j��  ]rD�  (j��  ]rE�  (j��  ]rF�  (h	h
e]rG�  (hh<e]rH�  (hhe]rI�  (j��  ]rJ�  (h	h
e]rK�  (hh�e]rL�  (hhe]rM�  (j��  ]rN�  (h	he]rO�  (hh�eeee]rP�  (hhee]rQ�  (h!]rR�  (h#h$e]rS�  (h	j�  e]rT�  (hh�e]rU�  (h)heeejC�  jC�  ]rV�  (j��  ]rW�  (j��  ]rX�  (j��  ]rY�  (h	h
e]rZ�  (hh<e]r[�  (hhe]r\�  (j��  ]r]�  (h	h
e]r^�  (hh�e]r_�  (hhe]r`�  (j��  ]ra�  (h	he]rb�  (hh�eeee]rc�  (hhee]rd�  (h!]re�  (h#h$e]rf�  (h	j�  e]rg�  (hh�e]rh�  (h)heeejV�  ]ri�  (j��  ]rj�  (j��  ]rk�  (j��  ]rl�  (h	h
e]rm�  (hh<e]rn�  (hhe]ro�  (j��  ]rp�  (h	h
e]rq�  (hh�e]rr�  (hhe]rs�  (j��  ]rt�  (h	he]ru�  (hh�eeee]rv�  (hhee]rw�  (h!]rx�  (h#h$e]ry�  (h	j�  e]rz�  (hh�e]r{�  (h)heeeji�  ]r|�  (j��  ]r}�  (j��  ]r~�  (j��  ]r�  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r  (hhee]r×  (h!]rė  (h#h$e]rŗ  (h	j�  e]rƗ  (hh�e]rǗ  (h)heeej��  j��  ]rȗ  (j��  ]rɗ  (j��  ]rʗ  (j��  ]r˗  (h	h
e]r̗  (hh<e]r͗  (hhe]rΗ  (j��  ]rϗ  (h	h
e]rЗ  (hh�e]rї  (hhe]rҗ  (j��  ]rӗ  (h	he]rԗ  (hh�eeee]r՗  (hhee]r֗  (h!]rח  (h#h$e]rؗ  (h	j�  e]rٗ  (hh�e]rڗ  (h)heeejȗ  jȗ  ]rۗ  (j��  ]rܗ  (j��  ]rݗ  (j��  ]rޗ  (h	h
e]rߗ  (hh<e]r��  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r �  (h)heeej�  j�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r	�  (hh�e]r
�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (X	   Next-Mover�  ]r �  (h	he]r!�  (hh�eeee]r"�  (hhee]r#�  (h!]r$�  (h#h$e]r%�  (h	j�  e]r&�  (hh<e]r'�  (h)heeej�  ]r(�  (j��  ]r)�  (j��  ]r*�  (j��  ]r+�  (h	h
e]r,�  (hh<e]r-�  (hhe]r.�  (j��  ]r/�  (h	h
e]r0�  (hh�e]r1�  (hhe]r2�  (j�  ]r3�  (h	he]r4�  (hh�eeee]r5�  (hhee]r6�  (h!]r7�  (h#h$e]r8�  (h	j�  e]r9�  (hh<e]r:�  (h)heeej(�  j(�  j(�  j(�  ]r;�  (j��  ]r<�  (j��  ]r=�  (j��  ]r>�  (h	h
e]r?�  (hh<e]r@�  (hhe]rA�  (j��  ]rB�  (h	h
e]rC�  (hh�e]rD�  (hhe]rE�  (j�  ]rF�  (h	he]rG�  (hh�eeee]rH�  (hhee]rI�  (h!]rJ�  (h#h$e]rK�  (h	he]rL�  (hh<e]rM�  (h)heee]rN�  (j��  ]rO�  (j��  ]rP�  (j��  ]rQ�  (h	h
e]rR�  (hh<e]rS�  (hhe]rT�  (j��  ]rU�  (h	h
e]rV�  (hh�e]rW�  (hhe]rX�  (j�  ]rY�  (h	he]rZ�  (hh�eeee]r[�  (hhee]r\�  (h!]r]�  (h#h$e]r^�  (h	he]r_�  (hh<e]r`�  (h)heeejN�  ]ra�  (j��  ]rb�  (j��  ]rc�  (j��  ]rd�  (h	h
e]re�  (hh<e]rf�  (hhe]rg�  (j��  ]rh�  (h	h
e]ri�  (hh�e]rj�  (hhe]rk�  (j�  ]rl�  (h	he]rm�  (hh�eeee]rn�  (hhee]ro�  (h!]rp�  (h#h$e]rq�  (h	h�e]rr�  (hh<e]rs�  (h)heeeja�  ja�  ja�  ]rt�  (j��  ]ru�  (j��  ]rv�  (j��  ]rw�  (h	h
e]rx�  (hh�e]ry�  (hhe]rz�  (j��  ]r{�  (h	h
e]r|�  (hh�e]r}�  (hhe]r~�  (j�  ]r�  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh<e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh<e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh<e]r��  (h)heeej��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh<e]r��  (h)heeej��  j��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r  (j��  ]rØ  (h	h
e]rĘ  (hh�e]rŘ  (hhe]rƘ  (j��  ]rǘ  (h	h
e]rȘ  (hh�e]rɘ  (hhe]rʘ  (j�  ]r˘  (h	he]r̘  (hh�eeee]r͘  (hhee]rΘ  (h!]rϘ  (h#h$e]rИ  (h	h�e]rј  (hh<e]rҘ  (h)heeej��  ]rӘ  (j��  ]rԘ  (j��  ]r՘  (j��  ]r֘  (h	h
e]rט  (hh�e]rؘ  (hhe]r٘  (j��  ]rژ  (h	h
e]rۘ  (hh�e]rܘ  (hhe]rݘ  (j�  ]rޘ  (h	he]rߘ  (hh�eeee]r��  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh<e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r��  (h!]r��  (h#h$e]r��  (h	he]r��  (hh<e]r��  (h)heeej�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r �  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r	�  (h	he]r
�  (hh<e]r�  (h)heeej��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh<e]r�  (h)heeej�  j�  j�  j�  j�  ]r�  (j��  ]r �  (j��  ]r!�  (j��  ]r"�  (h	h
e]r#�  (hh�e]r$�  (hhe]r%�  (j��  ]r&�  (h	h
e]r'�  (hh�e]r(�  (hhe]r)�  (j�  ]r*�  (h	he]r+�  (hh�eeee]r,�  (hhee]r-�  (h!]r.�  (h#h$e]r/�  (h	he]r0�  (hh�e]r1�  (h)heee]r2�  (j��  ]r3�  (j��  ]r4�  (j��  ]r5�  (h	h
e]r6�  (hh�e]r7�  (hhe]r8�  (j��  ]r9�  (h	h
e]r:�  (hh�e]r;�  (hhe]r<�  (j�  ]r=�  (h	he]r>�  (hh�eeee]r?�  (hhee]r@�  (h!]rA�  (h#h$e]rB�  (h	j�  e]rC�  (hh�e]rD�  (h)heeej2�  j2�  ]rE�  (j��  ]rF�  (j��  ]rG�  (j��  ]rH�  (h	h
e]rI�  (hh�e]rJ�  (hhe]rK�  (j��  ]rL�  (h	h
e]rM�  (hh�e]rN�  (hhe]rO�  (j�  ]rP�  (h	he]rQ�  (hh�eeee]rR�  (hhee]rS�  (h!]rT�  (h#h$e]rU�  (h	h�e]rV�  (hh�e]rW�  (h)heee]rX�  (j��  ]rY�  (j��  ]rZ�  (j��  ]r[�  (h	h
e]r\�  (hh�e]r]�  (hhe]r^�  (j��  ]r_�  (h	h
e]r`�  (hh�e]ra�  (hhe]rb�  (j�  ]rc�  (h	he]rd�  (hh�eeee]re�  (hhee]rf�  (h!]rg�  (h#h$e]rh�  (h	h�e]ri�  (hh�e]rj�  (h)heeejX�  jX�  ]rk�  (j��  ]rl�  (j��  ]rm�  (j��  ]rn�  (h	h
e]ro�  (hh�e]rp�  (hhe]rq�  (j��  ]rr�  (h	h
e]rs�  (hh<e]rt�  (hhe]ru�  (j�  ]rv�  (h	he]rw�  (hh�eeee]rx�  (hhee]ry�  (h!]rz�  (h#h$e]r{�  (h	h�e]r|�  (hh�e]r}�  (h)heeejk�  ]r~�  (j��  ]r�  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej~�  j~�  j~�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)h�eeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)h�eeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r  (h	he]rÙ  (hh�eeee]rę  (hhee]rř  (h!]rƙ  (h#h$e]rǙ  (h	j�  e]rș  (hh<e]rə  (h)h�eeej��  j��  ]rʙ  (j��  ]r˙  (j��  ]r̙  (j��  ]r͙  (h	h
e]rΙ  (hh�e]rϙ  (hhe]rЙ  (j��  ]rљ  (h	h
e]rҙ  (hh<e]rә  (hhe]rԙ  (j�  ]rՙ  (h	he]r֙  (hh�eeee]rי  (hhee]rؙ  (h!]rٙ  (h#h$e]rڙ  (h	j�  e]rۙ  (hh<e]rܙ  (h)h�eeejʙ  ]rݙ  (j��  ]rޙ  (j��  ]rߙ  (j��  ]r��  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r �  (h	j�  e]r�  (hh<e]r�  (h)heeej�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r	�  (j��  ]r
�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	j�  e]r�  (hh<e]r�  (h)heeej�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r �  (j�  ]r!�  (h	h�e]r"�  (hh�eeee]r#�  (hhee]r$�  (h!]r%�  (h#h$e]r&�  (h	j�  e]r'�  (hh<e]r(�  (h)heee]r)�  (j��  ]r*�  (j��  ]r+�  (j��  ]r,�  (h	h
e]r-�  (hh�e]r.�  (hhe]r/�  (j��  ]r0�  (h	h
e]r1�  (hh<e]r2�  (hhe]r3�  (j�  ]r4�  (h	he]r5�  (hh�eeee]r6�  (hhee]r7�  (h!]r8�  (h#h$e]r9�  (h	j�  e]r:�  (hh<e]r;�  (h)heee]r<�  (j��  ]r=�  (j��  ]r>�  (j��  ]r?�  (h	h
e]r@�  (hh�e]rA�  (hhe]rB�  (j��  ]rC�  (h	h
e]rD�  (hh<e]rE�  (hhe]rF�  (j�  ]rG�  (h	he]rH�  (hh�eeee]rI�  (hhee]rJ�  (h!]rK�  (h#h$e]rL�  (h	j�  e]rM�  (hh<e]rN�  (h)heeej<�  j<�  j<�  ]rO�  (j��  ]rP�  (j��  ]rQ�  (j��  ]rR�  (h	h
e]rS�  (hh�e]rT�  (hhe]rU�  (j��  ]rV�  (h	h
e]rW�  (hh<e]rX�  (hhe]rY�  (j�  ]rZ�  (h	he]r[�  (hh�eeee]r\�  (hhee]r]�  (h!]r^�  (h#h$e]r_�  (h	j�  e]r`�  (hh<e]ra�  (h)h�eee]rb�  (j��  ]rc�  (j��  ]rd�  (j��  ]re�  (h	h
e]rf�  (hh�e]rg�  (hhe]rh�  (j��  ]ri�  (h	h
e]rj�  (hh<e]rk�  (hhe]rl�  (j�  ]rm�  (h	he]rn�  (hh�eeee]ro�  (hhee]rp�  (h!]rq�  (h#h$e]rr�  (h	j�  e]rs�  (hh<e]rt�  (h)h�eee]ru�  (j��  ]rv�  (j��  ]rw�  (j��  ]rx�  (h	h
e]ry�  (hh�e]rz�  (hhe]r{�  (j��  ]r|�  (h	h
e]r}�  (hh�e]r~�  (hhe]r�  (j�  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)h�eee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)h�eee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)h�eeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh<e]r��  (h)h�eeej��  ]r��  (j��  ]r  (j��  ]rÚ  (j��  ]rĚ  (h	h
e]rŚ  (hh�e]rƚ  (hhe]rǚ  (j��  ]rȚ  (h	h
e]rɚ  (hh�e]rʚ  (hhe]r˚  (j�  ]r̚  (h	he]r͚  (hh�eeee]rΚ  (hhee]rϚ  (h!]rК  (h#h$e]rњ  (h	j�  e]rҚ  (hh<e]rӚ  (h)heeej��  j��  j��  j��  j��  j��  ]rԚ  (j��  ]r՚  (j��  ]r֚  (j��  ]rך  (h	h
e]rؚ  (hh�e]rٚ  (hhe]rښ  (j��  ]rۚ  (h	h
e]rܚ  (hh�e]rݚ  (hhe]rޚ  (j�  ]rߚ  (h	he]r��  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r �  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r	�  (h#h$e]r
�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  ]r �  (j��  ]r!�  (j��  ]r"�  (j��  ]r#�  (h	h
e]r$�  (hh�e]r%�  (hhe]r&�  (j��  ]r'�  (h	h
e]r(�  (hh<e]r)�  (hhe]r*�  (j�  ]r+�  (h	he]r,�  (hh�eeee]r-�  (hhee]r.�  (h!]r/�  (h#h$e]r0�  (h	h�e]r1�  (hh�e]r2�  (h)heeej �  ]r3�  (j��  ]r4�  (j��  ]r5�  (j��  ]r6�  (h	h
e]r7�  (hh�e]r8�  (hhe]r9�  (j��  ]r:�  (h	h
e]r;�  (hh<e]r<�  (hhe]r=�  (j�  ]r>�  (h	he]r?�  (hh�eeee]r@�  (hhee]rA�  (h!]rB�  (h#h$e]rC�  (h	h�e]rD�  (hh�e]rE�  (h)heeej3�  j3�  ]rF�  (j��  ]rG�  (j��  ]rH�  (j��  ]rI�  (h	h
e]rJ�  (hh�e]rK�  (hhe]rL�  (j��  ]rM�  (h	h
e]rN�  (hh<e]rO�  (hhe]rP�  (j�  ]rQ�  (h	he]rR�  (hh�eeee]rS�  (hhee]rT�  (h!]rU�  (h#h$e]rV�  (h	j�  e]rW�  (hh�e]rX�  (h)heee]rY�  (j��  ]rZ�  (j��  ]r[�  (j��  ]r\�  (h	h
e]r]�  (hh�e]r^�  (hhe]r_�  (j��  ]r`�  (h	h
e]ra�  (hh<e]rb�  (hhe]rc�  (j�  ]rd�  (h	he]re�  (hh�eeee]rf�  (hhee]rg�  (h!]rh�  (h#h$e]ri�  (h	he]rj�  (hh�e]rk�  (h)heeejY�  jY�  jY�  ]rl�  (j��  ]rm�  (j��  ]rn�  (j��  ]ro�  (h	h
e]rp�  (hh�e]rq�  (hhe]rr�  (j��  ]rs�  (h	h
e]rt�  (hh<e]ru�  (hhe]rv�  (j�  ]rw�  (h	h�e]rx�  (hh�eeee]ry�  (hhee]rz�  (h!]r{�  (h#h$e]r|�  (h	he]r}�  (hh�e]r~�  (h)heeejl�  jl�  jl�  ]r�  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)heeej�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r  (j�  ]rÛ  (h	h�e]rě  (hh�eeee]rś  (hhee]rƛ  (h!]rǛ  (h#h$e]rț  (h	h
e]rɛ  (hh�e]rʛ  (h)heee]r˛  (j��  ]r̛  (j��  ]r͛  (j��  ]rΛ  (h	h
e]rϛ  (hh�e]rЛ  (hhe]rћ  (j��  ]rқ  (h	h
e]rӛ  (hh�e]rԛ  (hhe]r՛  (j�  ]r֛  (h	h�e]rכ  (hh�eeee]r؛  (hhee]rٛ  (h!]rڛ  (h#h$e]rۛ  (h	h
e]rܛ  (hh�e]rݛ  (h)heeej˛  ]rޛ  (j��  ]rߛ  (j��  ]r��  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heeejޛ  jޛ  jޛ  jޛ  jޛ  jޛ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r �  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r	�  (hhe]r
�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)h�eeej�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r �  (hhe]r!�  (j�  ]r"�  (h	h�e]r#�  (hh�eeee]r$�  (hhee]r%�  (h!]r&�  (h#h$e]r'�  (h	h
e]r(�  (hh�e]r)�  (h)h�eee]r*�  (j��  ]r+�  (j��  ]r,�  (j��  ]r-�  (h	h
e]r.�  (hh<e]r/�  (hhe]r0�  (j��  ]r1�  (h	h
e]r2�  (hh�e]r3�  (hhe]r4�  (j�  ]r5�  (h	h�e]r6�  (hh�eeee]r7�  (hhee]r8�  (h!]r9�  (h#h$e]r:�  (h	j�  e]r;�  (hh�e]r<�  (h)h�eeej*�  j*�  j*�  j*�  ]r=�  (j��  ]r>�  (j��  ]r?�  (j��  ]r@�  (h	h
e]rA�  (hh<e]rB�  (hhe]rC�  (j��  ]rD�  (h	h
e]rE�  (hh�e]rF�  (hhe]rG�  (j�  ]rH�  (h	h�e]rI�  (hh�eeee]rJ�  (hhee]rK�  (h!]rL�  (h#h$e]rM�  (h	h
e]rN�  (hh�e]rO�  (h)h�eee]rP�  (j��  ]rQ�  (j��  ]rR�  (j��  ]rS�  (h	h
e]rT�  (hh<e]rU�  (hhe]rV�  (j��  ]rW�  (h	h
e]rX�  (hh�e]rY�  (hhe]rZ�  (j�  ]r[�  (h	h�e]r\�  (hh�eeee]r]�  (hhee]r^�  (h!]r_�  (h#h$e]r`�  (h	h
e]ra�  (hh�e]rb�  (h)heeejP�  jP�  ]rc�  (j��  ]rd�  (j��  ]re�  (j��  ]rf�  (h	h
e]rg�  (hh<e]rh�  (hhe]ri�  (j��  ]rj�  (h	h
e]rk�  (hh�e]rl�  (hhe]rm�  (j�  ]rn�  (h	h�e]ro�  (hh�eeee]rp�  (hhee]rq�  (h!]rr�  (h#h$e]rs�  (h	h
e]rt�  (hh�e]ru�  (h)heee]rv�  (j��  ]rw�  (j��  ]rx�  (j��  ]ry�  (h	h�e]rz�  (hh<e]r{�  (hhe]r|�  (j��  ]r}�  (h	h
e]r~�  (hh�e]r�  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heeejv�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r  (j��  ]rÜ  (j��  ]rĜ  (j��  ]rŜ  (h	h�e]rƜ  (hh<e]rǜ  (hhe]rȜ  (j��  ]rɜ  (h	h
e]rʜ  (hh<e]r˜  (hhe]r̜  (j�  ]r͜  (h	h�e]rΜ  (hh�eeee]rϜ  (hhee]rМ  (h!]rќ  (h#h$e]rҜ  (h	h�e]rӜ  (hh�e]rԜ  (h)heeej  ]r՜  (j��  ]r֜  (j��  ]rל  (j��  ]r؜  (h	h�e]rٜ  (hh<e]rڜ  (hhe]rۜ  (j��  ]rܜ  (h	h
e]rݜ  (hh<e]rޜ  (hhe]rߜ  (j�  ]r��  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r �  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r	�  (h!]r
�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heeej��  j��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r �  (h)heeej�  j�  ]r!�  (j��  ]r"�  (j��  ]r#�  (j��  ]r$�  (h	h�e]r%�  (hh<e]r&�  (hhe]r'�  (j��  ]r(�  (h	h�e]r)�  (hh<e]r*�  (hhe]r+�  (j�  ]r,�  (h	h�e]r-�  (hh�eeee]r.�  (hhee]r/�  (h!]r0�  (h#h$e]r1�  (h	h
e]r2�  (hh�e]r3�  (h)heee]r4�  (j��  ]r5�  (j��  ]r6�  (j��  ]r7�  (h	h�e]r8�  (hh<e]r9�  (hhe]r:�  (j��  ]r;�  (h	h�e]r<�  (hh<e]r=�  (hhe]r>�  (j�  ]r?�  (h	h�e]r@�  (hh�eeee]rA�  (hhee]rB�  (h!]rC�  (h#h$e]rD�  (h	h
e]rE�  (hh�e]rF�  (h)heee]rG�  (j��  ]rH�  (j��  ]rI�  (j��  ]rJ�  (h	h�e]rK�  (hh<e]rL�  (hhe]rM�  (j��  ]rN�  (h	h�e]rO�  (hh<e]rP�  (hhe]rQ�  (j�  ]rR�  (h	h�e]rS�  (hh�eeee]rT�  (hhee]rU�  (h!]rV�  (h#h$e]rW�  (h	h
e]rX�  (hh�e]rY�  (h)heee]rZ�  (j��  ]r[�  (j��  ]r\�  (j��  ]r]�  (h	h�e]r^�  (hh<e]r_�  (hhe]r`�  (j��  ]ra�  (h	h�e]rb�  (hh<e]rc�  (hhe]rd�  (j�  ]re�  (h	h�e]rf�  (hh�eeee]rg�  (hhee]rh�  (h!]ri�  (h#h$e]rj�  (h	h
e]rk�  (hh�e]rl�  (h)heee]rm�  (j��  ]rn�  (j��  ]ro�  (j��  ]rp�  (h	h�e]rq�  (hh<e]rr�  (hhe]rs�  (j��  ]rt�  (h	h�e]ru�  (hh<e]rv�  (hhe]rw�  (j�  ]rx�  (h	h�e]ry�  (hh�eeee]rz�  (hhee]r{�  (h!]r|�  (h#h$e]r}�  (h	h
e]r~�  (hh�e]r�  (h)heeejm�  jm�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h
e]r��  (hh<e]r��  (h)heeej��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r  (hhe]rÝ  (j�  ]rĝ  (h	h�e]rŝ  (hh�eeee]rƝ  (hhee]rǝ  (h!]rȝ  (h#h$e]rɝ  (h	h
e]rʝ  (hh�e]r˝  (h)heee]r̝  (j��  ]r͝  (j��  ]rΝ  (j��  ]rϝ  (h	h�e]rН  (hh<e]rѝ  (hhe]rҝ  (j��  ]rӝ  (h	h�e]rԝ  (hh<e]r՝  (hhe]r֝  (j�  ]rם  (h	h�e]r؝  (hh�eeee]rٝ  (hhee]rڝ  (h!]r۝  (h#h$e]rܝ  (h	h
e]rݝ  (hh�e]rޝ  (h)heeej̝  ]rߝ  (j��  ]r��  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heeejߝ  jߝ  ]r�  (j��  ]r�  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r �  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r	�  (hh<e]r
�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h
e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r �  (hh<e]r!�  (hhe]r"�  (j�  ]r#�  (h	h�e]r$�  (hh�eeee]r%�  (hhee]r&�  (h!]r'�  (h#h$e]r(�  (h	h
e]r)�  (hh�e]r*�  (h)heee]r+�  (j��  ]r,�  (j��  ]r-�  (j��  ]r.�  (h	h�e]r/�  (hh<e]r0�  (hhe]r1�  (j��  ]r2�  (h	h�e]r3�  (hh<e]r4�  (hhe]r5�  (j�  ]r6�  (h	h�e]r7�  (hh�eeee]r8�  (hhee]r9�  (h!]r:�  (h#h$e]r;�  (h	h
e]r<�  (hh�e]r=�  (h)heeej+�  ]r>�  (j��  ]r?�  (j��  ]r@�  (j��  ]rA�  (h	h�e]rB�  (hh<e]rC�  (hhe]rD�  (j��  ]rE�  (h	h
e]rF�  (hh<e]rG�  (hhe]rH�  (j�  ]rI�  (h	h�e]rJ�  (hh�eeee]rK�  (hhee]rL�  (h!]rM�  (h#h$e]rN�  (h	h
e]rO�  (hh�e]rP�  (h)heee]rQ�  (j��  ]rR�  (j��  ]rS�  (j��  ]rT�  (h	h�e]rU�  (hh<e]rV�  (hhe]rW�  (j��  ]rX�  (h	h
e]rY�  (hh<e]rZ�  (hhe]r[�  (j�  ]r\�  (h	h�e]r]�  (hh�eeee]r^�  (hhee]r_�  (h!]r`�  (h#h$e]ra�  (h	h
e]rb�  (hh<e]rc�  (h)heeejQ�  jQ�  ]rd�  (j��  ]re�  (j��  ]rf�  (j��  ]rg�  (h	h�e]rh�  (hh<e]ri�  (hhe]rj�  (j��  ]rk�  (h	h
e]rl�  (hh<e]rm�  (hhe]rn�  (j�  ]ro�  (h	h�e]rp�  (hh�eeee]rq�  (hhee]rr�  (h!]rs�  (h#h$e]rt�  (h	j�  e]ru�  (hh�e]rv�  (h)h�eeejd�  ]rw�  (j��  ]rx�  (j��  ]ry�  (j��  ]rz�  (h	h
e]r{�  (hh<e]r|�  (hhe]r}�  (j��  ]r~�  (h	h
e]r�  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)h�eee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)h�eeej��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r��  (h)h�eee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	j�  e]r��  (hh�e]r  (h)heeej��  j��  ]rÞ  (j��  ]rĞ  (j��  ]rŞ  (j��  ]rƞ  (h	h
e]rǞ  (hh�e]rȞ  (hhe]rɞ  (j��  ]rʞ  (h	h
e]r˞  (hh<e]r̞  (hhe]r͞  (j�  ]rΞ  (h	h�e]rϞ  (hh�eeee]rО  (hhee]rў  (h!]rҞ  (h#h$e]rӞ  (h	he]rԞ  (hh�e]r՞  (h)heeejÞ  ]r֞  (j��  ]rמ  (j��  ]r؞  (j��  ]rٞ  (h	h
e]rڞ  (hh�e]r۞  (hhe]rܞ  (j��  ]rݞ  (h	h
e]rޞ  (hh<e]rߞ  (hhe]r��  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	he]r�  (hh�e]r�  (h)heeej֞  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r �  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r	�  (hhee]r
�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  j��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r �  (hh�e]r!�  (h)heee]r"�  (j��  ]r#�  (j��  ]r$�  (j��  ]r%�  (h	h
e]r&�  (hh�e]r'�  (hhe]r(�  (j��  ]r)�  (h	h
e]r*�  (hh<e]r+�  (hhe]r,�  (j�  ]r-�  (h	h�e]r.�  (hh�eeee]r/�  (hhee]r0�  (h!]r1�  (h#h$e]r2�  (h	h�e]r3�  (hh�e]r4�  (h)heeej"�  ]r5�  (j��  ]r6�  (j��  ]r7�  (j��  ]r8�  (h	h
e]r9�  (hh�e]r:�  (hhe]r;�  (j��  ]r<�  (h	h
e]r=�  (hh<e]r>�  (hhe]r?�  (j�  ]r@�  (h	h�e]rA�  (hh�eeee]rB�  (hhee]rC�  (h!]rD�  (h#h$e]rE�  (h	h�e]rF�  (hh�e]rG�  (h)heeej5�  j5�  j5�  ]rH�  (j��  ]rI�  (j��  ]rJ�  (j��  ]rK�  (h	h
e]rL�  (hh�e]rM�  (hhe]rN�  (j��  ]rO�  (h	h
e]rP�  (hh<e]rQ�  (hhe]rR�  (j�  ]rS�  (h	h�e]rT�  (hh�eeee]rU�  (hhee]rV�  (h!]rW�  (h#h$e]rX�  (h	h�e]rY�  (hh�e]rZ�  (h)h�eee]r[�  (j��  ]r\�  (j��  ]r]�  (j��  ]r^�  (h	h
e]r_�  (hh�e]r`�  (hhe]ra�  (j��  ]rb�  (h	h
e]rc�  (hh<e]rd�  (hhe]re�  (j�  ]rf�  (h	h�e]rg�  (hh�eeee]rh�  (hhee]ri�  (h!]rj�  (h#h$e]rk�  (h	h�e]rl�  (hh�e]rm�  (h)h�eeej[�  j[�  j[�  ]rn�  (j��  ]ro�  (j��  ]rp�  (j��  ]rq�  (h	h
e]rr�  (hh�e]rs�  (hhe]rt�  (j��  ]ru�  (h	h
e]rv�  (hh<e]rw�  (hhe]rx�  (j�  ]ry�  (h	h�e]rz�  (hh�eeee]r{�  (hhee]r|�  (h!]r}�  (h#h$e]r~�  (h	h�e]r�  (hh�e]r��  (h)h�eee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (X	   Next-Mover��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)h�eeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)h�eeej��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)h�eee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r  (h	h
e]rß  (hh<e]rğ  (hhe]rş  (j��  ]rƟ  (h	he]rǟ  (hh�eeee]rȟ  (hhee]rɟ  (h!]rʟ  (h#h$e]r˟  (h	h�e]r̟  (hh�e]r͟  (h)h�eee]rΟ  (j��  ]rϟ  (j��  ]rП  (j��  ]rџ  (h	h
e]rҟ  (hh�e]rӟ  (hhe]rԟ  (j��  ]r՟  (h	h
e]r֟  (hh<e]rן  (hhe]r؟  (j��  ]rٟ  (h	he]rڟ  (hh�eeee]r۟  (hhee]rܟ  (h!]rݟ  (h#h$e]rޟ  (h	h�e]rߟ  (hh�e]r��  (h)h�eeejΟ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)h�eee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	he]r �  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)h�eeej��  ]r�  (j��  ]r�  (j��  ]r	�  (j��  ]r
�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	he]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)h�eeej�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r �  (j��  ]r!�  (h	h
e]r"�  (hh<e]r#�  (hhe]r$�  (j��  ]r%�  (h	he]r&�  (hh�eeee]r'�  (hhee]r(�  (h!]r)�  (h#h$e]r*�  (h	h�e]r+�  (hh�e]r,�  (h)h�eee]r-�  (j��  ]r.�  (j��  ]r/�  (j��  ]r0�  (h	h
e]r1�  (hh�e]r2�  (hhe]r3�  (j��  ]r4�  (h	h
e]r5�  (hh<e]r6�  (hhe]r7�  (X	   Next-Mover8�  ]r9�  (h	h�e]r:�  (hh�eeee]r;�  (hhee]r<�  (h!]r=�  (h#h$e]r>�  (h	h�e]r?�  (hh�e]r@�  (h)h�eee]rA�  (j��  ]rB�  (j��  ]rC�  (j��  ]rD�  (h	h
e]rE�  (hh�e]rF�  (hhe]rG�  (j��  ]rH�  (h	h
e]rI�  (hh<e]rJ�  (hhe]rK�  (j8�  ]rL�  (h	h�e]rM�  (hh�eeee]rN�  (hhee]rO�  (h!]rP�  (h#h$e]rQ�  (h	h�e]rR�  (hh�e]rS�  (h)h�eeejA�  ]rT�  (j��  ]rU�  (j��  ]rV�  (j��  ]rW�  (h	h
e]rX�  (hh�e]rY�  (hhe]rZ�  (j��  ]r[�  (h	h
e]r\�  (hh<e]r]�  (hhe]r^�  (j8�  ]r_�  (h	h�e]r`�  (hh�eeee]ra�  (hhee]rb�  (h!]rc�  (h#h$e]rd�  (h	h�e]re�  (hh�e]rf�  (h)heeejT�  jT�  jT�  ]rg�  (j��  ]rh�  (j��  ]ri�  (j��  ]rj�  (h	h
e]rk�  (hh�e]rl�  (hhe]rm�  (j��  ]rn�  (h	h
e]ro�  (hh<e]rp�  (hhe]rq�  (j8�  ]rr�  (h	h�e]rs�  (hh�eeee]rt�  (hhee]ru�  (h!]rv�  (h#h$e]rw�  (h	h�e]rx�  (hh�e]ry�  (h)heeejg�  ]rz�  (j��  ]r{�  (j��  ]r|�  (j��  ]r}�  (h	h
e]r~�  (hh�e]r�  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeejz�  jz�  jz�  jz�  jz�  jz�  jz�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r   (h#h$e]rà  (h	h�e]rĠ  (hh�e]rŠ  (h)heeej��  ]rƠ  (j��  ]rǠ  (j��  ]rȠ  (j��  ]rɠ  (h	h
e]rʠ  (hh�e]rˠ  (hhe]r̠  (j��  ]r͠  (h	h
e]rΠ  (hh�e]rϠ  (hhe]rР  (j8�  ]rѠ  (h	h�e]rҠ  (hh�eeee]rӠ  (hhee]rԠ  (h!]rՠ  (h#h$e]r֠  (h	h�e]rנ  (hh�e]rؠ  (h)heeejƠ  jƠ  jƠ  jƠ  ]r٠  (j��  ]rڠ  (j��  ]r۠  (j��  ]rܠ  (h	h
e]rݠ  (hh�e]rޠ  (hhe]rߠ  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej٠  j٠  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  ]r��  (j��  ]r �  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r	�  (j8�  ]r
�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej��  j��  j��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r �  (h!]r!�  (h#h$e]r"�  (h	h�e]r#�  (hh�e]r$�  (h)heeej�  j�  j�  j�  ]r%�  (j��  ]r&�  (j��  ]r'�  (j��  ]r(�  (h	h
e]r)�  (hh<e]r*�  (hhe]r+�  (j��  ]r,�  (h	h
e]r-�  (hh�e]r.�  (hhe]r/�  (j8�  ]r0�  (h	h�e]r1�  (hh�eeee]r2�  (hhee]r3�  (h!]r4�  (h#h$e]r5�  (h	h�e]r6�  (hh�e]r7�  (h)heeej%�  j%�  j%�  j%�  j%�  j%�  j%�  j%�  j%�  j%�  j%�  j%�  j%�  ]r8�  (j��  ]r9�  (j��  ]r:�  (j��  ]r;�  (h	h
e]r<�  (hh<e]r=�  (hhe]r>�  (j��  ]r?�  (h	h
e]r@�  (hh�e]rA�  (hhe]rB�  (j8�  ]rC�  (h	h�e]rD�  (hh�eeee]rE�  (hhee]rF�  (h!]rG�  (h#h$e]rH�  (h	h�e]rI�  (hh�e]rJ�  (h)heeej8�  ]rK�  (j��  ]rL�  (j��  ]rM�  (j��  ]rN�  (h	h
e]rO�  (hh<e]rP�  (hhe]rQ�  (j��  ]rR�  (h	h
e]rS�  (hh�e]rT�  (hhe]rU�  (j8�  ]rV�  (h	h�e]rW�  (hh�eeee]rX�  (hhee]rY�  (h!]rZ�  (h#h$e]r[�  (h	h�e]r\�  (hh�e]r]�  (h)heeejK�  jK�  ]r^�  (j��  ]r_�  (j��  ]r`�  (j��  ]ra�  (h	h
e]rb�  (hh<e]rc�  (hhe]rd�  (j��  ]re�  (h	h
e]rf�  (hh�e]rg�  (hhe]rh�  (j8�  ]ri�  (h	h�e]rj�  (hh�eeee]rk�  (hhee]rl�  (h!]rm�  (h#h$e]rn�  (h	h�e]ro�  (hh�e]rp�  (h)heeej^�  ]rq�  (j��  ]rr�  (j��  ]rs�  (j��  ]rt�  (h	h
e]ru�  (hh<e]rv�  (hhe]rw�  (j��  ]rx�  (h	h
e]ry�  (hh�e]rz�  (hhe]r{�  (j8�  ]r|�  (h	h�e]r}�  (hh�eeee]r~�  (hhee]r�  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r¡  (hhe]rá  (j��  ]rġ  (h	h
e]rš  (hh�e]rơ  (hhe]rǡ  (j8�  ]rȡ  (h	h�e]rɡ  (hh�eeee]rʡ  (hhee]rˡ  (h!]r̡  (h#h$e]r͡  (h	h�e]rΡ  (hh�e]rϡ  (h)heee]rС  (j��  ]rѡ  (j��  ]rҡ  (j��  ]rӡ  (h	h
e]rԡ  (hh<e]rա  (hhe]r֡  (j��  ]rס  (h	h
e]rء  (hh�e]r١  (hhe]rڡ  (j8�  ]rۡ  (h	h�e]rܡ  (hh�eeee]rݡ  (hhee]rޡ  (h!]rߡ  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejС  jС  jС  jС  jС  jС  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r �  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r	�  (j��  ]r
�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej	�  j	�  j	�  j	�  j	�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r �  (hh<e]r!�  (hhe]r"�  (j��  ]r#�  (h	h
e]r$�  (hh�e]r%�  (hhe]r&�  (j8�  ]r'�  (h	h�e]r(�  (hh�eeee]r)�  (hhee]r*�  (h!]r+�  (h#h$e]r,�  (h	h�e]r-�  (hh�e]r.�  (h)heeej�  j�  ]r/�  (j��  ]r0�  (j��  ]r1�  (j��  ]r2�  (h	h
e]r3�  (hh<e]r4�  (hhe]r5�  (j��  ]r6�  (h	h
e]r7�  (hh�e]r8�  (hhe]r9�  (j8�  ]r:�  (h	h�e]r;�  (hh�eeee]r<�  (hhee]r=�  (h!]r>�  (h#h$e]r?�  (h	h�e]r@�  (hh�e]rA�  (h)heee]rB�  (j��  ]rC�  (j��  ]rD�  (j��  ]rE�  (h	h
e]rF�  (hh<e]rG�  (hhe]rH�  (j��  ]rI�  (h	h
e]rJ�  (hh�e]rK�  (hhe]rL�  (j8�  ]rM�  (h	h�e]rN�  (hh�eeee]rO�  (hhee]rP�  (h!]rQ�  (h#h$e]rR�  (h	h�e]rS�  (hh�e]rT�  (h)heeejB�  jB�  ]rU�  (j��  ]rV�  (j��  ]rW�  (j��  ]rX�  (h	h
e]rY�  (hh<e]rZ�  (hhe]r[�  (j��  ]r\�  (h	h
e]r]�  (hh�e]r^�  (hhe]r_�  (j8�  ]r`�  (h	h�e]ra�  (hh�eeee]rb�  (hhee]rc�  (h!]rd�  (h#h$e]re�  (h	h�e]rf�  (hh�e]rg�  (h)heeejU�  jU�  jU�  jU�  jU�  jU�  ]rh�  (j��  ]ri�  (j��  ]rj�  (j��  ]rk�  (h	h
e]rl�  (hh<e]rm�  (hhe]rn�  (j��  ]ro�  (h	h
e]rp�  (hh�e]rq�  (hhe]rr�  (j8�  ]rs�  (h	h�e]rt�  (hh�eeee]ru�  (hhee]rv�  (h!]rw�  (h#h$e]rx�  (h	h�e]ry�  (hh�e]rz�  (h)heeejh�  ]r{�  (j��  ]r|�  (j��  ]r}�  (j��  ]r~�  (h	h
e]r�  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej{�  j{�  j{�  j{�  j{�  j{�  j{�  j{�  j{�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r¢  (h!]râ  (h#h$e]rĢ  (h	h�e]rŢ  (hh�e]rƢ  (h)heee]rǢ  (j��  ]rȢ  (j��  ]rɢ  (j��  ]rʢ  (h	h
e]rˢ  (hh<e]r̢  (hhe]r͢  (j��  ]r΢  (h	h
e]rϢ  (hh�e]rТ  (hhe]rѢ  (j8�  ]rҢ  (h	h�e]rӢ  (hh�eeee]rԢ  (hhee]rբ  (h!]r֢  (h#h$e]rע  (h	h�e]rآ  (hh�e]r٢  (h)heeejǢ  jǢ  jǢ  jǢ  jǢ  jǢ  jǢ  jǢ  jǢ  jǢ  jǢ  ]rڢ  (j��  ]rۢ  (j��  ]rܢ  (j��  ]rݢ  (h	h
e]rޢ  (hh<e]rߢ  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejڢ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  ]r �  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r	�  (hhe]r
�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r �  (hhee]r!�  (h!]r"�  (h#h$e]r#�  (h	h�e]r$�  (hh�e]r%�  (h)heeej�  j�  ]r&�  (j��  ]r'�  (j��  ]r(�  (j��  ]r)�  (h	h�e]r*�  (hh<e]r+�  (hhe]r,�  (j��  ]r-�  (h	h
e]r.�  (hh<e]r/�  (hhe]r0�  (j8�  ]r1�  (h	h�e]r2�  (hh�eeee]r3�  (hhee]r4�  (h!]r5�  (h#h$e]r6�  (h	h�e]r7�  (hh�e]r8�  (h)heee]r9�  (j��  ]r:�  (j��  ]r;�  (j��  ]r<�  (h	h�e]r=�  (hh<e]r>�  (hhe]r?�  (j��  ]r@�  (h	h
e]rA�  (hh<e]rB�  (hhe]rC�  (j8�  ]rD�  (h	h�e]rE�  (hh�eeee]rF�  (hhee]rG�  (h!]rH�  (h#h$e]rI�  (h	h�e]rJ�  (hh�e]rK�  (h)heeej9�  j9�  j9�  j9�  j9�  j9�  j9�  j9�  j9�  j9�  j9�  ]rL�  (j��  ]rM�  (j��  ]rN�  (j��  ]rO�  (h	h�e]rP�  (hh<e]rQ�  (hhe]rR�  (j��  ]rS�  (h	h
e]rT�  (hh<e]rU�  (hhe]rV�  (j8�  ]rW�  (h	h�e]rX�  (hh�eeee]rY�  (hhee]rZ�  (h!]r[�  (h#h$e]r\�  (h	h�e]r]�  (hh�e]r^�  (h)heeejL�  ]r_�  (j��  ]r`�  (j��  ]ra�  (j��  ]rb�  (h	h�e]rc�  (hh<e]rd�  (hhe]re�  (j��  ]rf�  (h	h
e]rg�  (hh<e]rh�  (hhe]ri�  (j8�  ]rj�  (h	h�e]rk�  (hh�eeee]rl�  (hhee]rm�  (h!]rn�  (h#h$e]ro�  (h	h�e]rp�  (hh�e]rq�  (h)heee]rr�  (j��  ]rs�  (j��  ]rt�  (j��  ]ru�  (h	h�e]rv�  (hh<e]rw�  (hhe]rx�  (j��  ]ry�  (h	h
e]rz�  (hh<e]r{�  (hhe]r|�  (j8�  ]r}�  (h	h�e]r~�  (hh�eeee]r�  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeejr�  jr�  jr�  jr�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r£  (hh<e]rã  (hhe]rģ  (j��  ]rţ  (h	h
e]rƣ  (hh<e]rǣ  (hhe]rȣ  (j8�  ]rɣ  (h	h�e]rʣ  (hh�eeee]rˣ  (hhee]ṛ  (h!]rͣ  (h#h$e]rΣ  (h	h�e]rϣ  (hh�e]rУ  (h)heeej��  ]rѣ  (j��  ]rң  (j��  ]rӣ  (j��  ]rԣ  (h	h�e]rգ  (hh<e]r֣  (hhe]rף  (j��  ]rأ  (h	h
e]r٣  (hh<e]rڣ  (hhe]rۣ  (j8�  ]rܣ  (h	h�e]rݣ  (hh�eeee]rޣ  (hhee]rߣ  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejѣ  jѣ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r �  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r	�  (h)heeej��  j��  ]r
�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej
�  j
�  j
�  j
�  j
�  j
�  j
�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r �  (h	h�e]r!�  (hh<e]r"�  (hhe]r#�  (j��  ]r$�  (h	h
e]r%�  (hh�e]r&�  (hhe]r'�  (j8�  ]r(�  (h	h�e]r)�  (hh�eeee]r*�  (hhee]r+�  (h!]r,�  (h#h$e]r-�  (h	h�e]r.�  (hh�e]r/�  (h)heeej�  j�  ]r0�  (j��  ]r1�  (j��  ]r2�  (j��  ]r3�  (h	h�e]r4�  (hh<e]r5�  (hhe]r6�  (j��  ]r7�  (h	h
e]r8�  (hh�e]r9�  (hhe]r:�  (j8�  ]r;�  (h	h�e]r<�  (hh�eeee]r=�  (hhee]r>�  (h!]r?�  (h#h$e]r@�  (h	h�e]rA�  (hh�e]rB�  (h)heeej0�  j0�  j0�  j0�  j0�  j0�  j0�  j0�  j0�  j0�  ]rC�  (j��  ]rD�  (j��  ]rE�  (j��  ]rF�  (h	h�e]rG�  (hh<e]rH�  (hhe]rI�  (j��  ]rJ�  (h	h
e]rK�  (hh�e]rL�  (hhe]rM�  (j8�  ]rN�  (h	h�e]rO�  (hh�eeee]rP�  (hhee]rQ�  (h!]rR�  (h#h$e]rS�  (h	h�e]rT�  (hh�e]rU�  (h)heeejC�  jC�  jC�  jC�  ]rV�  (j��  ]rW�  (j��  ]rX�  (j��  ]rY�  (h	h�e]rZ�  (hh<e]r[�  (hhe]r\�  (j��  ]r]�  (h	h
e]r^�  (hh�e]r_�  (hhe]r`�  (j8�  ]ra�  (h	h�e]rb�  (hh�eeee]rc�  (hhee]rd�  (h!]re�  (h#h$e]rf�  (h	h�e]rg�  (hh�e]rh�  (h)heeejV�  jV�  jV�  jV�  ]ri�  (j��  ]rj�  (j��  ]rk�  (j��  ]rl�  (h	h�e]rm�  (hh<e]rn�  (hhe]ro�  (j��  ]rp�  (h	h
e]rq�  (hh<e]rr�  (hhe]rs�  (j8�  ]rt�  (h	h�e]ru�  (hh�eeee]rv�  (hhee]rw�  (h!]rx�  (h#h$e]ry�  (h	h�e]rz�  (hh�e]r{�  (h)heeeji�  ji�  ji�  ]r|�  (j��  ]r}�  (j��  ]r~�  (j��  ]r�  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej|�  j|�  j|�  j|�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r¤  (hhee]rä  (h!]rĤ  (h#h$e]rŤ  (h	h�e]rƤ  (hh�e]rǤ  (h)heee]rȤ  (j��  ]rɤ  (j��  ]rʤ  (j��  ]rˤ  (h	h�e]r̤  (hh<e]rͤ  (hhe]rΤ  (j��  ]rϤ  (h	h
e]rФ  (hh<e]rѤ  (hhe]rҤ  (j8�  ]rӤ  (h	h�e]rԤ  (hh�eeee]rդ  (hhee]r֤  (h!]rפ  (h#h$e]rؤ  (h	h�e]r٤  (hh�e]rڤ  (h)heeejȤ  jȤ  jȤ  jȤ  jȤ  jȤ  ]rۤ  (j��  ]rܤ  (j��  ]rݤ  (j��  ]rޤ  (h	h�e]rߤ  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejۤ  jۤ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r �  (h)heeej�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r	�  (hh<e]r
�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeee(j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r �  (hh�eeee]r!�  (hhee]r"�  (h!]r#�  (h#h$e]r$�  (h	h�e]r%�  (hh�e]r&�  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r'�  (j��  ]r(�  (j��  ]r)�  (j��  ]r*�  (h	h�e]r+�  (hh<e]r,�  (hhe]r-�  (j��  ]r.�  (h	h�e]r/�  (hh<e]r0�  (hhe]r1�  (j8�  ]r2�  (h	h�e]r3�  (hh�eeee]r4�  (hhee]r5�  (h!]r6�  (h#h$e]r7�  (h	h�e]r8�  (hh�e]r9�  (h)heeej'�  j'�  j'�  j'�  ]r:�  (j��  ]r;�  (j��  ]r<�  (j��  ]r=�  (h	h�e]r>�  (hh<e]r?�  (hhe]r@�  (j��  ]rA�  (h	h�e]rB�  (hh<e]rC�  (hhe]rD�  (j8�  ]rE�  (h	h�e]rF�  (hh�eeee]rG�  (hhee]rH�  (h!]rI�  (h#h$e]rJ�  (h	h�e]rK�  (hh�e]rL�  (h)heeej:�  ]rM�  (j��  ]rN�  (j��  ]rO�  (j��  ]rP�  (h	h�e]rQ�  (hh<e]rR�  (hhe]rS�  (j��  ]rT�  (h	h�e]rU�  (hh<e]rV�  (hhe]rW�  (j8�  ]rX�  (h	h�e]rY�  (hh�eeee]rZ�  (hhee]r[�  (h!]r\�  (h#h$e]r]�  (h	h�e]r^�  (hh�e]r_�  (h)heee]r`�  (j��  ]ra�  (j��  ]rb�  (j��  ]rc�  (h	h�e]rd�  (hh<e]re�  (hhe]rf�  (j��  ]rg�  (h	h�e]rh�  (hh<e]ri�  (hhe]rj�  (j8�  ]rk�  (h	h�e]rl�  (hh�eeee]rm�  (hhee]rn�  (h!]ro�  (h#h$e]rp�  (h	h�e]rq�  (hh�e]rr�  (h)heeej`�  j`�  j`�  j`�  j`�  j`�  ]rs�  (j��  ]rt�  (j��  ]ru�  (j��  ]rv�  (h	h�e]rw�  (hh<e]rx�  (hhe]ry�  (j��  ]rz�  (h	h�e]r{�  (hh<e]r|�  (hhe]r}�  (j8�  ]r~�  (h	h�e]r�  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeejs�  js�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r¥  (h	h�e]rå  (hh<e]rĥ  (hhe]rť  (j��  ]rƥ  (h	h�e]rǥ  (hh<e]rȥ  (hhe]rɥ  (j8�  ]rʥ  (h	h�e]r˥  (hh�eeee]r̥  (hhee]rͥ  (h!]rΥ  (h#h$e]rϥ  (h	h�e]rХ  (hh�e]rѥ  (h)heee]rҥ  (j��  ]rӥ  (j��  ]rԥ  (j��  ]rե  (h	h�e]r֥  (hh<e]rץ  (hhe]rإ  (j��  ]r٥  (h	h�e]rڥ  (hh<e]rۥ  (hhe]rܥ  (j8�  ]rݥ  (h	h�e]rޥ  (hh�eeee]rߥ  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejҥ  jҥ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r �  (hh<e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r	�  (hh�e]r
�  (h)heeej��  j��  j��  j��  j��  j��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j8�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (j��  ]r�  (j��  ]r �  (j��  ]r!�  (h	h�e]r"�  (hh<e]r#�  (hhe]r$�  (j��  ]r%�  (h	h�e]r&�  (hh<e]r'�  (hhe]r(�  (j8�  ]r)�  (h	h�e]r*�  (hh�eeee]r+�  (hhee]r,�  (h!]r-�  (h#h$e]r.�  (h	h�e]r/�  (hh�e]r0�  (h)heee]r1�  (j��  ]r2�  (j��  ]r3�  (j��  ]r4�  (h	h�e]r5�  (hh<e]r6�  (hhe]r7�  (j��  ]r8�  (h	h�e]r9�  (hh<e]r:�  (hhe]r;�  (j8�  ]r<�  (h	h�e]r=�  (hh�eeee]r>�  (hhee]r?�  (h!]r@�  (h#h$e]rA�  (h	h�e]rB�  (hh�e]rC�  (h)heeej1�  j1�  j1�  j1�  j1�  j1�  j1�  j1�  ]rD�  (j��  ]rE�  (j��  ]rF�  (j��  ]rG�  (h	h
e]rH�  (hh<e]rI�  (hhe]rJ�  (j��  ]rK�  (h	h�e]rL�  (hh<e]rM�  (hhe]rN�  (j8�  ]rO�  (h	h�e]rP�  (hh�eeee]rQ�  (hhee]rR�  (h!]rS�  (h#h$e]rT�  (h	h�e]rU�  (hh�e]rV�  (h)heeejD�  ]rW�  (j��  ]rX�  (j��  ]rY�  (j��  ]rZ�  (h	h
e]r[�  (hh<e]r\�  (hhe]r]�  (j��  ]r^�  (h	h�e]r_�  (hh<e]r`�  (hhe]ra�  (j8�  ]rb�  (h	h�e]rc�  (hh�eeee]rd�  (hhee]re�  (h!]rf�  (h#h$e]rg�  (h	h�e]rh�  (hh�e]ri�  (h)heeejW�  jW�  jW�  ]rj�  (j��  ]rk�  (j��  ]rl�  (j��  ]rm�  (h	h�e]rn�  (hh<e]ro�  (hhe]rp�  (j��  ]rq�  (h	h�e]rr�  (hh<e]rs�  (hhe]rt�  (j8�  ]ru�  (h	h�e]rv�  (hh�eeee]rw�  (hhee]rx�  (h!]ry�  (h#h$e]rz�  (h	h�e]r{�  (hh�e]r|�  (h)heee]r}�  (j��  ]r~�  (j��  ]r�  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j8�  ]r��  (h	h�e]r¦  (hh�eeee]ræ  (hhee]rĦ  (h!]rŦ  (h#h$e]rƦ  (h	h�e]rǦ  (hh�e]rȦ  (h)heeej��  j��  j��  j��  ]rɦ  (j��  ]rʦ  (j��  ]r˦  (j��  ]r̦  (h	h�e]rͦ  (hh<e]rΦ  (hhe]rϦ  (j��  ]rЦ  (h	h
e]rѦ  (hh<e]rҦ  (hhe]rӦ  (j8�  ]rԦ  (h	h�e]rզ  (hh�eeee]r֦  (hhee]rצ  (h!]rئ  (h#h$e]r٦  (h	h�e]rڦ  (hh�e]rۦ  (h)heee]rܦ  (j��  ]rݦ  (j��  ]rަ  (j��  ]rߦ  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (X	   Next-Mover�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r �  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r	�  (j��  ]r
�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r �  (j�  ]r!�  (h	h�e]r"�  (hh�eeee]r#�  (hhee]r$�  (h!]r%�  (h#h$e]r&�  (h	h�e]r'�  (hh�e]r(�  (h)heeej�  ]r)�  (j��  ]r*�  (j��  ]r+�  (j��  ]r,�  (h	h�e]r-�  (hh<e]r.�  (hhe]r/�  (j��  ]r0�  (h	h
e]r1�  (hh<e]r2�  (hhe]r3�  (j�  ]r4�  (h	h�e]r5�  (hh�eeee]r6�  (hhee]r7�  (h!]r8�  (h#h$e]r9�  (h	h�e]r:�  (hh�e]r;�  (h)heee]r<�  (j��  ]r=�  (j��  ]r>�  (j��  ]r?�  (h	h�e]r@�  (hh<e]rA�  (hhe]rB�  (j��  ]rC�  (h	h
e]rD�  (hh<e]rE�  (hhe]rF�  (j�  ]rG�  (h	h�e]rH�  (hh�eeee]rI�  (hhee]rJ�  (h!]rK�  (h#h$e]rL�  (h	h�e]rM�  (hh�e]rN�  (h)heeej<�  j<�  j<�  j<�  j<�  j<�  j<�  j<�  j<�  ]rO�  (j��  ]rP�  (j��  ]rQ�  (j��  ]rR�  (h	h�e]rS�  (hh<e]rT�  (hhe]rU�  (j��  ]rV�  (h	h
e]rW�  (hh<e]rX�  (hhe]rY�  (j�  ]rZ�  (h	h�e]r[�  (hh�eeee]r\�  (hhee]r]�  (h!]r^�  (h#h$e]r_�  (h	h�e]r`�  (hh�e]ra�  (h)heeejO�  ]rb�  (j��  ]rc�  (j��  ]rd�  (j��  ]re�  (h	h�e]rf�  (hh<e]rg�  (hhe]rh�  (j��  ]ri�  (h	h
e]rj�  (hh<e]rk�  (hhe]rl�  (j�  ]rm�  (h	h�e]rn�  (hh�eeee]ro�  (hhee]rp�  (h!]rq�  (h#h$e]rr�  (h	h�e]rs�  (hh�e]rt�  (h)heeejb�  jb�  jb�  jb�  ]ru�  (j��  ]rv�  (j��  ]rw�  (j��  ]rx�  (h	h�e]ry�  (hh<e]rz�  (hhe]r{�  (j��  ]r|�  (h	h
e]r}�  (hh<e]r~�  (hhe]r�  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeeju�  ju�  ju�  ju�  ju�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r§  (j��  ]rç  (j��  ]rħ  (h	h�e]rŧ  (hh<e]rƧ  (hhe]rǧ  (j��  ]rȧ  (h	h�e]rɧ  (hh<e]rʧ  (hhe]r˧  (j�  ]ŗ  (h	h�e]rͧ  (hh�eeee]rΧ  (hhee]rϧ  (h!]rЧ  (h#h$e]rѧ  (h	h�e]rҧ  (hh�e]rӧ  (h)heee]rԧ  (j��  ]rէ  (j��  ]r֧  (j��  ]rק  (h	h�e]rا  (hh<e]r٧  (hhe]rڧ  (j��  ]rۧ  (h	h�e]rܧ  (hh<e]rݧ  (hhe]rާ  (j�  ]rߧ  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejԧ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r �  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r	�  (h#h$e]r
�  (h	h�e]r�  (hh�e]r�  (h)heeej��  j��  j��  j��  j��  j��  j��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r �  (j��  ]r!�  (j��  ]r"�  (j��  ]r#�  (h	h�e]r$�  (hh<e]r%�  (hhe]r&�  (j��  ]r'�  (h	h
e]r(�  (hh<e]r)�  (hhe]r*�  (j�  ]r+�  (h	h�e]r,�  (hh�eeee]r-�  (hhee]r.�  (h!]r/�  (h#h$e]r0�  (h	h�e]r1�  (hh�e]r2�  (h)heeej �  ]r3�  (j��  ]r4�  (j��  ]r5�  (j��  ]r6�  (h	h
e]r7�  (hh<e]r8�  (hhe]r9�  (j��  ]r:�  (h	h
e]r;�  (hh<e]r<�  (hhe]r=�  (j�  ]r>�  (h	h�e]r?�  (hh�eeee]r@�  (hhee]rA�  (h!]rB�  (h#h$e]rC�  (h	h�e]rD�  (hh�e]rE�  (h)heeej3�  ]rF�  (j��  ]rG�  (j��  ]rH�  (j��  ]rI�  (h	h
e]rJ�  (hh<e]rK�  (hhe]rL�  (j��  ]rM�  (h	h
e]rN�  (hh<e]rO�  (hhe]rP�  (j�  ]rQ�  (h	h�e]rR�  (hh�eeee]rS�  (hhee]rT�  (h!]rU�  (h#h$e]rV�  (h	h�e]rW�  (hh�e]rX�  (h)heeejF�  jF�  ]rY�  (j��  ]rZ�  (j��  ]r[�  (j��  ]r\�  (h	h
e]r]�  (hh<e]r^�  (hhe]r_�  (j��  ]r`�  (h	h
e]ra�  (hh<e]rb�  (hhe]rc�  (j�  ]rd�  (h	h�e]re�  (hh�eeee]rf�  (hhee]rg�  (h!]rh�  (h#h$e]ri�  (h	h�e]rj�  (hh�e]rk�  (h)heeejY�  jY�  ]rl�  (j��  ]rm�  (j��  ]rn�  (j��  ]ro�  (h	h
e]rp�  (hh<e]rq�  (hhe]rr�  (j��  ]rs�  (h	h
e]rt�  (hh<e]ru�  (hhe]rv�  (j�  ]rw�  (h	h�e]rx�  (hh�eeee]ry�  (hhee]rz�  (h!]r{�  (h#h$e]r|�  (h	h�e]r}�  (hh�e]r~�  (h)heee]r�  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r¨  (j�  ]rè  (h	h�e]rĨ  (hh�eeee]rŨ  (hhee]rƨ  (h!]rǨ  (h#h$e]rȨ  (h	h�e]rɨ  (hh�e]rʨ  (h)heee]r˨  (j��  ]r̨  (j��  ]rͨ  (j��  ]rΨ  (h	h
e]rϨ  (hh<e]rШ  (hhe]rѨ  (j��  ]rҨ  (h	h�e]rӨ  (hh<e]rԨ  (hhe]rը  (j�  ]r֨  (h	h�e]rר  (hh�eeee]rب  (hhee]r٨  (h!]rڨ  (h#h$e]rۨ  (h	h�e]rܨ  (hh�e]rݨ  (h)heee]rި  (j��  ]rߨ  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejި  jި  jި  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r �  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r	�  (hhe]r
�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r �  (hhe]r!�  (j�  ]r"�  (h	h�e]r#�  (hh�eeee]r$�  (hhee]r%�  (h!]r&�  (h#h$e]r'�  (h	h�e]r(�  (hh�e]r)�  (h)heee]r*�  (j��  ]r+�  (j��  ]r,�  (j��  ]r-�  (h	h
e]r.�  (hh<e]r/�  (hhe]r0�  (j��  ]r1�  (h	h�e]r2�  (hh<e]r3�  (hhe]r4�  (j�  ]r5�  (h	h�e]r6�  (hh�eeee]r7�  (hhee]r8�  (h!]r9�  (h#h$e]r:�  (h	h�e]r;�  (hh�e]r<�  (h)heeej*�  j*�  j*�  j*�  j*�  j*�  j*�  j*�  j*�  j*�  ]r=�  (j��  ]r>�  (j��  ]r?�  (j��  ]r@�  (h	h
e]rA�  (hh<e]rB�  (hhe]rC�  (j��  ]rD�  (h	h�e]rE�  (hh<e]rF�  (hhe]rG�  (j�  ]rH�  (h	h�e]rI�  (hh�eeee]rJ�  (hhee]rK�  (h!]rL�  (h#h$e]rM�  (h	h�e]rN�  (hh�e]rO�  (h)heeej=�  j=�  j=�  ]rP�  (j��  ]rQ�  (j��  ]rR�  (j��  ]rS�  (h	h
e]rT�  (hh<e]rU�  (hhe]rV�  (j��  ]rW�  (h	h�e]rX�  (hh<e]rY�  (hhe]rZ�  (j�  ]r[�  (h	h�e]r\�  (hh�eeee]r]�  (hhee]r^�  (h!]r_�  (h#h$e]r`�  (h	h�e]ra�  (hh�e]rb�  (h)heee]rc�  (j��  ]rd�  (j��  ]re�  (j��  ]rf�  (h	h
e]rg�  (hh<e]rh�  (hhe]ri�  (j��  ]rj�  (h	h�e]rk�  (hh<e]rl�  (hhe]rm�  (j�  ]rn�  (h	h�e]ro�  (hh�eeee]rp�  (hhee]rq�  (h!]rr�  (h#h$e]rs�  (h	h�e]rt�  (hh�e]ru�  (h)heeejc�  jc�  ]rv�  (j��  ]rw�  (j��  ]rx�  (j��  ]ry�  (h	h
e]rz�  (hh<e]r{�  (hhe]r|�  (j��  ]r}�  (h	h�e]r~�  (hh<e]r�  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeejv�  jv�  jv�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  ]r©  (j��  ]ré  (j��  ]rĩ  (j��  ]rũ  (h	h�e]rƩ  (hh<e]rǩ  (hhe]rȩ  (j��  ]rɩ  (h	h�e]rʩ  (hh<e]r˩  (hhe]r̩  (j�  ]rͩ  (h	h�e]rΩ  (hh�eeee]rϩ  (hhee]rЩ  (h!]rѩ  (h#h$e]rҩ  (h	h�e]rө  (hh�e]rԩ  (h)heee]rթ  (j��  ]r֩  (j��  ]rש  (j��  ]rة  (h	h�e]r٩  (hh<e]rک  (hhe]r۩  (j��  ]rܩ  (h	h�e]rݩ  (hh<e]rީ  (hhe]rߩ  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejթ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r �  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r	�  (h!]r
�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  j��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r �  (h)heeej�  ]r!�  (j��  ]r"�  (j��  ]r#�  (j��  ]r$�  (h	h
e]r%�  (hh<e]r&�  (hhe]r'�  (j��  ]r(�  (h	h�e]r)�  (hh<e]r*�  (hhe]r+�  (j�  ]r,�  (h	h�e]r-�  (hh�eeee]r.�  (hhee]r/�  (h!]r0�  (h#h$e]r1�  (h	h�e]r2�  (hh�e]r3�  (h)heee]r4�  (j��  ]r5�  (j��  ]r6�  (j��  ]r7�  (h	h
e]r8�  (hh<e]r9�  (hhe]r:�  (j��  ]r;�  (h	h�e]r<�  (hh<e]r=�  (hhe]r>�  (j�  ]r?�  (h	h�e]r@�  (hh�eeee]rA�  (hhee]rB�  (h!]rC�  (h#h$e]rD�  (h	h�e]rE�  (hh�e]rF�  (h)heeej4�  j4�  j4�  j4�  ]rG�  (j��  ]rH�  (j��  ]rI�  (j��  ]rJ�  (h	h
e]rK�  (hh<e]rL�  (hhe]rM�  (j��  ]rN�  (h	h�e]rO�  (hh<e]rP�  (hhe]rQ�  (j�  ]rR�  (h	h�e]rS�  (hh�eeee]rT�  (hhee]rU�  (h!]rV�  (h#h$e]rW�  (h	h�e]rX�  (hh�e]rY�  (h)heeejG�  jG�  jG�  jG�  jG�  jG�  jG�  ]rZ�  (j��  ]r[�  (j��  ]r\�  (j��  ]r]�  (h	h
e]r^�  (hh�e]r_�  (hhe]r`�  (j��  ]ra�  (h	h�e]rb�  (hh<e]rc�  (hhe]rd�  (j�  ]re�  (h	h�e]rf�  (hh�eeee]rg�  (hhee]rh�  (h!]ri�  (h#h$e]rj�  (h	h�e]rk�  (hh�e]rl�  (h)heeejZ�  jZ�  jZ�  jZ�  jZ�  jZ�  jZ�  ]rm�  (j��  ]rn�  (j��  ]ro�  (j��  ]rp�  (h	h
e]rq�  (hh�e]rr�  (hhe]rs�  (j��  ]rt�  (h	h
e]ru�  (hh<e]rv�  (hhe]rw�  (j�  ]rx�  (h	h�e]ry�  (hh�eeee]rz�  (hhee]r{�  (h!]r|�  (h#h$e]r}�  (h	h�e]r~�  (hh�e]r�  (h)heeejm�  jm�  jm�  jm�  jm�  jm�  jm�  jm�  jm�  jm�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]rª  (hhe]rê  (j�  ]rĪ  (h	h�e]rŪ  (hh�eeee]rƪ  (hhee]rǪ  (h!]rȪ  (h#h$e]rɪ  (h	h�e]rʪ  (hh�e]r˪  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  ]r̪  (j��  ]rͪ  (j��  ]rΪ  (j��  ]rϪ  (h	h
e]rЪ  (hh<e]rѪ  (hhe]rҪ  (j��  ]rӪ  (h	h
e]rԪ  (hh<e]rժ  (hhe]r֪  (j�  ]rת  (h	h�e]rت  (hh�eeee]r٪  (hhee]rڪ  (h!]r۪  (h#h$e]rܪ  (h	h�e]rݪ  (hh�e]rު  (h)heeej̪  ]rߪ  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejߪ  ]r�  (j��  ]r�  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r �  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r	�  (hh<e]r
�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r �  (hh<e]r!�  (hhe]r"�  (j�  ]r#�  (h	h�e]r$�  (hh�eeee]r%�  (hhee]r&�  (h!]r'�  (h#h$e]r(�  (h	h�e]r)�  (hh�e]r*�  (h)heee]r+�  (j��  ]r,�  (j��  ]r-�  (j��  ]r.�  (h	h
e]r/�  (hh�e]r0�  (hhe]r1�  (j��  ]r2�  (h	h
e]r3�  (hh<e]r4�  (hhe]r5�  (j�  ]r6�  (h	h�e]r7�  (hh�eeee]r8�  (hhee]r9�  (h!]r:�  (h#h$e]r;�  (h	h�e]r<�  (hh�e]r=�  (h)heee]r>�  (j��  ]r?�  (j��  ]r@�  (j��  ]rA�  (h	h
e]rB�  (hh�e]rC�  (hhe]rD�  (j��  ]rE�  (h	h
e]rF�  (hh<e]rG�  (hhe]rH�  (j�  ]rI�  (h	h�e]rJ�  (hh�eeee]rK�  (hhee]rL�  (h!]rM�  (h#h$e]rN�  (h	h�e]rO�  (hh�e]rP�  (h)heeej>�  j>�  j>�  ]rQ�  (j��  ]rR�  (j��  ]rS�  (j��  ]rT�  (h	h
e]rU�  (hh�e]rV�  (hhe]rW�  (j��  ]rX�  (h	h
e]rY�  (hh<e]rZ�  (hhe]r[�  (j�  ]r\�  (h	h�e]r]�  (hh�eeee]r^�  (hhee]r_�  (h!]r`�  (h#h$e]ra�  (h	h�e]rb�  (hh�e]rc�  (h)heee]rd�  (j��  ]re�  (j��  ]rf�  (j��  ]rg�  (h	h
e]rh�  (hh�e]ri�  (hhe]rj�  (j��  ]rk�  (h	h
e]rl�  (hh<e]rm�  (hhe]rn�  (j�  ]ro�  (h	h�e]rp�  (hh�eeee]rq�  (hhee]rr�  (h!]rs�  (h#h$e]rt�  (h	h�e]ru�  (hh�e]rv�  (h)heeejd�  jd�  ]rw�  (j��  ]rx�  (j��  ]ry�  (j��  ]rz�  (h	h
e]r{�  (hh�e]r|�  (hhe]r}�  (j��  ]r~�  (h	h
e]r�  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r«  (h)heeej��  j��  j��  ]rë  (j��  ]rī  (j��  ]rū  (j��  ]rƫ  (h	h
e]rǫ  (hh<e]rȫ  (hhe]rɫ  (j��  ]rʫ  (h	h
e]r˫  (hh<e]r̫  (hhe]rͫ  (j�  ]rΫ  (h	h�e]rϫ  (hh�eeee]rЫ  (hhee]rѫ  (h!]rҫ  (h#h$e]rӫ  (h	h�e]rԫ  (hh�e]rի  (h)heeejë  ]r֫  (j��  ]r׫  (j��  ]rث  (j��  ]r٫  (h	h
e]rګ  (hh<e]r۫  (hhe]rܫ  (j��  ]rݫ  (h	h
e]rޫ  (hh<e]r߫  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  j�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r �  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r	�  (hhee]r
�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej��  j��  j��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r �  (hh�e]r!�  (h)heeej�  ]r"�  (j��  ]r#�  (j��  ]r$�  (j��  ]r%�  (h	h
e]r&�  (hh<e]r'�  (hhe]r(�  (j��  ]r)�  (h	h�e]r*�  (hh<e]r+�  (hhe]r,�  (j�  ]r-�  (h	h�e]r.�  (hh�eeee]r/�  (hhee]r0�  (h!]r1�  (h#h$e]r2�  (h	h�e]r3�  (hh�e]r4�  (h)heee]r5�  (j��  ]r6�  (j��  ]r7�  (j��  ]r8�  (h	h
e]r9�  (hh<e]r:�  (hhe]r;�  (j��  ]r<�  (h	h�e]r=�  (hh<e]r>�  (hhe]r?�  (j�  ]r@�  (h	h�e]rA�  (hh�eeee]rB�  (hhee]rC�  (h!]rD�  (h#h$e]rE�  (h	h�e]rF�  (hh�e]rG�  (h)heeej5�  j5�  j5�  ]rH�  (j��  ]rI�  (j��  ]rJ�  (j��  ]rK�  (h	h
e]rL�  (hh<e]rM�  (hhe]rN�  (j��  ]rO�  (h	h�e]rP�  (hh<e]rQ�  (hhe]rR�  (j�  ]rS�  (h	h�e]rT�  (hh�eeee]rU�  (hhee]rV�  (h!]rW�  (h#h$e]rX�  (h	h�e]rY�  (hh�e]rZ�  (h)heeejH�  jH�  jH�  jH�  jH�  jH�  jH�  ]r[�  (j��  ]r\�  (j��  ]r]�  (j��  ]r^�  (h	h
e]r_�  (hh<e]r`�  (hhe]ra�  (j��  ]rb�  (h	h�e]rc�  (hh<e]rd�  (hhe]re�  (j�  ]rf�  (h	h�e]rg�  (hh�eeee]rh�  (hhee]ri�  (h!]rj�  (h#h$e]rk�  (h	h�e]rl�  (hh�e]rm�  (h)heeej[�  ]rn�  (j��  ]ro�  (j��  ]rp�  (j��  ]rq�  (h	h
e]rr�  (hh<e]rs�  (hhe]rt�  (j��  ]ru�  (h	h�e]rv�  (hh<e]rw�  (hhe]rx�  (j�  ]ry�  (h	h�e]rz�  (hh�eeee]r{�  (hhee]r|�  (h!]r}�  (h#h$e]r~�  (h	h�e]r�  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r¬  (hh<e]rì  (hhe]rĬ  (j�  ]rŬ  (h	h�e]rƬ  (hh�eeee]rǬ  (hhee]rȬ  (h!]rɬ  (h#h$e]rʬ  (h	h�e]rˬ  (hh�e]r̬  (h)heee]rͬ  (j��  ]rά  (j��  ]rϬ  (j��  ]rЬ  (h	h�e]rѬ  (hh<e]rҬ  (hhe]rӬ  (j��  ]rԬ  (h	h
e]rլ  (hh<e]r֬  (hhe]r׬  (j�  ]rج  (h	h�e]r٬  (hh�eeee]rڬ  (hhee]r۬  (h!]rܬ  (h#h$e]rݬ  (h	h�e]rެ  (hh�e]r߬  (h)heeejͬ  jͬ  jͬ  jͬ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r �  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r	�  (h	h
e]r
�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r �  (h	h
e]r!�  (hh<e]r"�  (hhe]r#�  (j�  ]r$�  (h	h�e]r%�  (hh�eeee]r&�  (hhee]r'�  (h!]r(�  (h#h$e]r)�  (h	h�e]r*�  (hh�e]r+�  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  j�  ]r,�  (j��  ]r-�  (j��  ]r.�  (j��  ]r/�  (h	h
e]r0�  (hh<e]r1�  (hhe]r2�  (j��  ]r3�  (h	h
e]r4�  (hh<e]r5�  (hhe]r6�  (j�  ]r7�  (h	h�e]r8�  (hh�eeee]r9�  (hhee]r:�  (h!]r;�  (h#h$e]r<�  (h	h�e]r=�  (hh�e]r>�  (h)heeej,�  ]r?�  (j��  ]r@�  (j��  ]rA�  (j��  ]rB�  (h	h
e]rC�  (hh<e]rD�  (hhe]rE�  (j��  ]rF�  (h	h
e]rG�  (hh<e]rH�  (hhe]rI�  (j�  ]rJ�  (h	h�e]rK�  (hh�eeee]rL�  (hhee]rM�  (h!]rN�  (h#h$e]rO�  (h	h�e]rP�  (hh�e]rQ�  (h)heee]rR�  (j��  ]rS�  (j��  ]rT�  (j��  ]rU�  (h	h
e]rV�  (hh<e]rW�  (hhe]rX�  (j��  ]rY�  (h	h
e]rZ�  (hh<e]r[�  (hhe]r\�  (j�  ]r]�  (h	h�e]r^�  (hh�eeee]r_�  (hhee]r`�  (h!]ra�  (h#h$e]rb�  (h	h�e]rc�  (hh�e]rd�  (h)heeejR�  jR�  ]re�  (j��  ]rf�  (j��  ]rg�  (j��  ]rh�  (h	h
e]ri�  (hh<e]rj�  (hhe]rk�  (j��  ]rl�  (h	h
e]rm�  (hh<e]rn�  (hhe]ro�  (j�  ]rp�  (h	h�e]rq�  (hh�eeee]rr�  (hhee]rs�  (h!]rt�  (h#h$e]ru�  (h	h�e]rv�  (hh�e]rw�  (h)heeeje�  je�  je�  ]rx�  (j��  ]ry�  (j��  ]rz�  (j��  ]r{�  (h	h
e]r|�  (hh<e]r}�  (hhe]r~�  (j��  ]r�  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r­  (hh�e]rí  (h)heee]rĭ  (j��  ]rŭ  (j��  ]rƭ  (j��  ]rǭ  (h	h
e]rȭ  (hh<e]rɭ  (hhe]rʭ  (j��  ]r˭  (h	h
e]r̭  (hh<e]rͭ  (hhe]rέ  (X	   Next-Moverϭ  ]rЭ  (h	h�e]rѭ  (hh�eeee]rҭ  (hhee]rӭ  (h!]rԭ  (h#h$e]rխ  (h	h�e]r֭  (hh�e]r׭  (h)heee]rح  (j��  ]r٭  (j��  ]rڭ  (j��  ]rۭ  (h	h
e]rܭ  (hh<e]rݭ  (hhe]rޭ  (j��  ]r߭  (h	h
e]r�  (hh<e]r�  (hhe]r�  (jϭ  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejح  jح  jح  jح  jح  jح  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r��  (hhe]r��  (jϭ  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r �  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (jϭ  ]r	�  (h	h�e]r
�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej��  j��  j��  j��  j��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (jϭ  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r �  (h#h$e]r!�  (h	h�e]r"�  (hh�e]r#�  (h)heeej�  ]r$�  (j��  ]r%�  (j��  ]r&�  (j��  ]r'�  (h	h
e]r(�  (hh<e]r)�  (hhe]r*�  (j��  ]r+�  (h	h�e]r,�  (hh<e]r-�  (hhe]r.�  (X	   Next-Mover/�  ]r0�  (h	h�e]r1�  (hh�eeee]r2�  (hhee]r3�  (h!]r4�  (h#h$e]r5�  (h	h�e]r6�  (hh�e]r7�  (h)heee]r8�  (j��  ]r9�  (j��  ]r:�  (j��  ]r;�  (h	h
e]r<�  (hh<e]r=�  (hhe]r>�  (j��  ]r?�  (h	h�e]r@�  (hh<e]rA�  (hhe]rB�  (j/�  ]rC�  (h	h�e]rD�  (hh�eeee]rE�  (hhee]rF�  (h!]rG�  (h#h$e]rH�  (h	h�e]rI�  (hh�e]rJ�  (h)heeej8�  ]rK�  (j��  ]rL�  (j��  ]rM�  (j��  ]rN�  (h	h
e]rO�  (hh<e]rP�  (hhe]rQ�  (j��  ]rR�  (h	h
e]rS�  (hh<e]rT�  (hhe]rU�  (j/�  ]rV�  (h	h�e]rW�  (hh�eeee]rX�  (hhee]rY�  (h!]rZ�  (h#h$e]r[�  (h	h�e]r\�  (hh�e]r]�  (h)heee]r^�  (j��  ]r_�  (j��  ]r`�  (j��  ]ra�  (h	h
e]rb�  (hh<e]rc�  (hhe]rd�  (j��  ]re�  (h	h�e]rf�  (hh<e]rg�  (hhe]rh�  (j/�  ]ri�  (h	h�e]rj�  (hh�eeee]rk�  (hhee]rl�  (h!]rm�  (h#h$e]rn�  (h	h�e]ro�  (hh�e]rp�  (h)heeej^�  ]rq�  (j��  ]rr�  (j��  ]rs�  (j��  ]rt�  (h	h
e]ru�  (hh<e]rv�  (hhe]rw�  (j��  ]rx�  (h	h�e]ry�  (hh<e]rz�  (hhe]r{�  (j/�  ]r|�  (h	h�e]r}�  (hh�eeee]r~�  (hhee]r�  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r®  (hhe]rî  (j��  ]rĮ  (h	h�e]rŮ  (hh<e]rƮ  (hhe]rǮ  (j/�  ]rȮ  (h	h�e]rɮ  (hh�eeee]rʮ  (hhee]rˮ  (h!]r̮  (h#h$e]rͮ  (h	h�e]rή  (hh�e]rϮ  (h)heeej��  j��  j��  ]rЮ  (j��  ]rѮ  (j��  ]rҮ  (j��  ]rӮ  (h	h�e]rԮ  (hh<e]rծ  (hhe]r֮  (j��  ]r׮  (h	h�e]rخ  (hh<e]rٮ  (hhe]rڮ  (j/�  ]rۮ  (h	h�e]rܮ  (hh�eeee]rݮ  (hhee]rޮ  (h!]r߮  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejЮ  jЮ  jЮ  jЮ  jЮ  jЮ  jЮ  jЮ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j/�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r �  (j/�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej��  j��  j��  ]r	�  (j��  ]r
�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j/�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej	�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r �  (hh<e]r!�  (hhe]r"�  (j��  ]r#�  (h	h�e]r$�  (hh<e]r%�  (hhe]r&�  (j/�  ]r'�  (h	h�e]r(�  (hh�eeee]r)�  (hhee]r*�  (h!]r+�  (h#h$e]r,�  (h	h�e]r-�  (hh�e]r.�  (h)heeej�  j�  j�  ]r/�  (j��  ]r0�  (j��  ]r1�  (j��  ]r2�  (h	h�e]r3�  (hh<e]r4�  (hhe]r5�  (j��  ]r6�  (h	h�e]r7�  (hh<e]r8�  (hhe]r9�  (j/�  ]r:�  (h	h�e]r;�  (hh�eeee]r<�  (hhee]r=�  (h!]r>�  (h#h$e]r?�  (h	h�e]r@�  (hh�e]rA�  (h)heee]rB�  (j��  ]rC�  (j��  ]rD�  (j��  ]rE�  (h	h�e]rF�  (hh<e]rG�  (hhe]rH�  (j��  ]rI�  (h	h�e]rJ�  (hh<e]rK�  (hhe]rL�  (j/�  ]rM�  (h	h�e]rN�  (hh�eeee]rO�  (hhee]rP�  (h!]rQ�  (h#h$e]rR�  (h	h�e]rS�  (hh�e]rT�  (h)heeejB�  jB�  jB�  jB�  jB�  ]rU�  (j��  ]rV�  (j��  ]rW�  (j��  ]rX�  (h	h�e]rY�  (hh<e]rZ�  (hhe]r[�  (j��  ]r\�  (h	h�e]r]�  (hh<e]r^�  (hhe]r_�  (j/�  ]r`�  (h	h�e]ra�  (hh�eeee]rb�  (hhee]rc�  (h!]rd�  (h#h$e]re�  (h	h�e]rf�  (hh�e]rg�  (h)heeejU�  ]rh�  (j��  ]ri�  (j��  ]rj�  (j��  ]rk�  (h	h�e]rl�  (hh<e]rm�  (hhe]rn�  (j��  ]ro�  (h	h�e]rp�  (hh<e]rq�  (hhe]rr�  (j/�  ]rs�  (h	h�e]rt�  (hh�eeee]ru�  (hhee]rv�  (h!]rw�  (h#h$e]rx�  (h	h�e]ry�  (hh�e]rz�  (h)heeejh�  jh�  jh�  jh�  jh�  jh�  ]r{�  (j��  ]r|�  (j��  ]r}�  (j��  ]r~�  (h	h�e]r�  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej{�  j{�  j{�  j{�  j{�  j{�  j{�  j{�  j{�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r¯  (h!]rï  (h#h$e]rį  (h	h�e]rů  (hh�e]rƯ  (h)heeej��  ]rǯ  (j��  ]rȯ  (j��  ]rɯ  (j��  ]rʯ  (h	h�e]r˯  (hh<e]r̯  (hhe]rͯ  (j��  ]rί  (h	h�e]rϯ  (hh<e]rЯ  (hhe]rѯ  (j/�  ]rү  (h	h�e]rӯ  (hh�eeee]rԯ  (hhee]rկ  (h!]r֯  (h#h$e]rׯ  (h	h�e]rد  (hh�e]rٯ  (h)heeejǯ  jǯ  jǯ  jǯ  jǯ  jǯ  jǯ  jǯ  ]rگ  (j��  ]rۯ  (j��  ]rܯ  (j��  ]rݯ  (h	h�e]rޯ  (hh<e]r߯  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j/�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejگ  jگ  jگ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  ]r �  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r	�  (hhe]r
�  (j/�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej �  j �  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j/�  ]r�  (h	h�e]r�  (hh�eeee]r �  (hhee]r!�  (h!]r"�  (h#h$e]r#�  (h	h�e]r$�  (hh�e]r%�  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  j�  ]r&�  (j��  ]r'�  (j��  ]r(�  (j��  ]r)�  (h	h�e]r*�  (hh<e]r+�  (hhe]r,�  (j��  ]r-�  (h	h�e]r.�  (hh<e]r/�  (hhe]r0�  (j/�  ]r1�  (h	h�e]r2�  (hh�eeee]r3�  (hhee]r4�  (h!]r5�  (h#h$e]r6�  (h	h�e]r7�  (hh�e]r8�  (h)heeej&�  ]r9�  (j��  ]r:�  (j��  ]r;�  (j��  ]r<�  (h	h�e]r=�  (hh<e]r>�  (hhe]r?�  (j��  ]r@�  (h	h�e]rA�  (hh<e]rB�  (hhe]rC�  (j/�  ]rD�  (h	h�e]rE�  (hh�eeee]rF�  (hhee]rG�  (h!]rH�  (h#h$e]rI�  (h	h�e]rJ�  (hh�e]rK�  (h)heeej9�  j9�  ]rL�  (j��  ]rM�  (j��  ]rN�  (j��  ]rO�  (h	h�e]rP�  (hh<e]rQ�  (hhe]rR�  (j��  ]rS�  (h	h
e]rT�  (hh<e]rU�  (hhe]rV�  (j/�  ]rW�  (h	h�e]rX�  (hh�eeee]rY�  (hhee]rZ�  (h!]r[�  (h#h$e]r\�  (h	h�e]r]�  (hh�e]r^�  (h)heeejL�  jL�  jL�  ]r_�  (j��  ]r`�  (j��  ]ra�  (j��  ]rb�  (h	h�e]rc�  (hh<e]rd�  (hhe]re�  (j��  ]rf�  (h	h
e]rg�  (hh<e]rh�  (hhe]ri�  (j/�  ]rj�  (h	h�e]rk�  (hh�eeee]rl�  (hhee]rm�  (h!]rn�  (h#h$e]ro�  (h	h�e]rp�  (hh�e]rq�  (h)heeej_�  ]rr�  (j��  ]rs�  (j��  ]rt�  (j��  ]ru�  (h	h�e]rv�  (hh<e]rw�  (hhe]rx�  (j��  ]ry�  (h	h
e]rz�  (hh<e]r{�  (hhe]r|�  (j/�  ]r}�  (h	h�e]r~�  (hh�eeee]r�  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeejr�  jr�  jr�  jr�  jr�  jr�  jr�  jr�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r°  (hh<e]rð  (hhe]rİ  (j��  ]rŰ  (h	h
e]rư  (hh<e]rǰ  (hhe]rȰ  (j/�  ]rɰ  (h	h�e]rʰ  (hh�eeee]r˰  (hhee]r̰  (h!]rͰ  (h#h$e]rΰ  (h	h�e]rϰ  (hh�e]rа  (h)heee]rѰ  (j��  ]rҰ  (j��  ]rӰ  (j��  ]r԰  (h	h�e]rհ  (hh<e]rְ  (hhe]rװ  (j��  ]rذ  (h	h
e]rٰ  (hh<e]rڰ  (hhe]r۰  (j/�  ]rܰ  (h	h�e]rݰ  (hh�eeee]rް  (hhee]r߰  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j/�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r �  (hhe]r�  (j/�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r	�  (h)heeej��  j��  j��  ]r
�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j/�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej
�  j
�  j
�  j
�  j
�  j
�  j
�  j
�  j
�  j
�  j
�  j
�  j
�  j
�  j
�  j
�  j
�  j
�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r �  (h	h�e]r!�  (hh<e]r"�  (hhe]r#�  (j��  ]r$�  (h	h
e]r%�  (hh<e]r&�  (hhe]r'�  (j/�  ]r(�  (h	h�e]r)�  (hh�eeee]r*�  (hhee]r+�  (h!]r,�  (h#h$e]r-�  (h	h�e]r.�  (hh�e]r/�  (h)heeej�  j�  j�  j�  j�  j�  j�  ]r0�  (j��  ]r1�  (j��  ]r2�  (j��  ]r3�  (h	h�e]r4�  (hh<e]r5�  (hhe]r6�  (j��  ]r7�  (h	h
e]r8�  (hh<e]r9�  (hhe]r:�  (j/�  ]r;�  (h	h�e]r<�  (hh�eeee]r=�  (hhee]r>�  (h!]r?�  (h#h$e]r@�  (h	h�e]rA�  (hh�e]rB�  (h)heeej0�  j0�  j0�  j0�  j0�  j0�  j0�  ]rC�  (j��  ]rD�  (j��  ]rE�  (j��  ]rF�  (h	h�e]rG�  (hh<e]rH�  (hhe]rI�  (j��  ]rJ�  (h	h
e]rK�  (hh<e]rL�  (hhe]rM�  (j/�  ]rN�  (h	h�e]rO�  (hh�eeee]rP�  (hhee]rQ�  (h!]rR�  (h#h$e]rS�  (h	h�e]rT�  (hh�e]rU�  (h)heeejC�  jC�  jC�  jC�  jC�  jC�  jC�  jC�  jC�  jC�  ]rV�  (j��  ]rW�  (j��  ]rX�  (j��  ]rY�  (h	h�e]rZ�  (hh<e]r[�  (hhe]r\�  (j��  ]r]�  (h	h
e]r^�  (hh<e]r_�  (hhe]r`�  (j/�  ]ra�  (h	h�e]rb�  (hh�eeee]rc�  (hhee]rd�  (h!]re�  (h#h$e]rf�  (h	h�e]rg�  (hh�e]rh�  (h)heeejV�  jV�  jV�  jV�  jV�  jV�  jV�  jV�  jV�  jV�  jV�  jV�  jV�  ]ri�  (j��  ]rj�  (j��  ]rk�  (j��  ]rl�  (h	h�e]rm�  (hh<e]rn�  (hhe]ro�  (j��  ]rp�  (h	h
e]rq�  (hh�e]rr�  (hhe]rs�  (j/�  ]rt�  (h	h�e]ru�  (hh�eeee]rv�  (hhee]rw�  (h!]rx�  (h#h$e]ry�  (h	h�e]rz�  (hh�e]r{�  (h)heeeji�  ji�  ji�  ji�  ji�  ji�  ji�  ji�  ]r|�  (j��  ]r}�  (j��  ]r~�  (j��  ]r�  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej|�  j|�  j|�  j|�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j/�  ]r��  (h	h�e]r��  (hh�eeee]r±  (hhee]rñ  (h!]rı  (h#h$e]rű  (h	h�e]rƱ  (hh�e]rǱ  (h)heeej��  j��  j��  j��  j��  ]rȱ  (j��  ]rɱ  (j��  ]rʱ  (j��  ]r˱  (h	h�e]ṟ  (hh<e]rͱ  (hhe]rα  (j��  ]rϱ  (h	h
e]rб  (hh�e]rѱ  (hhe]rұ  (j/�  ]rӱ  (h	h�e]rԱ  (hh�eeee]rձ  (hhee]rֱ  (h!]rױ  (h#h$e]rر  (h	h�e]rٱ  (hh�e]rڱ  (h)heeejȱ  jȱ  jȱ  ]r۱  (j��  ]rܱ  (j��  ]rݱ  (j��  ]rޱ  (h	h�e]r߱  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (X	   Next-Mover�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r �  (hh�e]r�  (h)heeej�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r	�  (h	h
e]r
�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j�  ]r �  (h	h�e]r!�  (hh�eeee]r"�  (hhee]r#�  (h!]r$�  (h#h$e]r%�  (h	h�e]r&�  (hh�e]r'�  (h)heeej�  ]r(�  (j��  ]r)�  (j��  ]r*�  (j��  ]r+�  (h	h�e]r,�  (hh<e]r-�  (hhe]r.�  (j��  ]r/�  (h	h
e]r0�  (hh�e]r1�  (hhe]r2�  (j�  ]r3�  (h	h�e]r4�  (hh�eeee]r5�  (hhee]r6�  (h!]r7�  (h#h$e]r8�  (h	h�e]r9�  (hh�e]r:�  (h)heee]r;�  (j��  ]r<�  (j��  ]r=�  (j��  ]r>�  (h	h�e]r?�  (hh<e]r@�  (hhe]rA�  (j��  ]rB�  (h	h
e]rC�  (hh�e]rD�  (hhe]rE�  (j�  ]rF�  (h	h�e]rG�  (hh�eeee]rH�  (hhee]rI�  (h!]rJ�  (h#h$e]rK�  (h	h�e]rL�  (hh�e]rM�  (h)heee]rN�  (j��  ]rO�  (j��  ]rP�  (j��  ]rQ�  (h	h�e]rR�  (hh<e]rS�  (hhe]rT�  (j��  ]rU�  (h	h
e]rV�  (hh�e]rW�  (hhe]rX�  (j�  ]rY�  (h	h�e]rZ�  (hh�eeee]r[�  (hhee]r\�  (h!]r]�  (h#h$e]r^�  (h	h�e]r_�  (hh�e]r`�  (h)heeejN�  ]ra�  (j��  ]rb�  (j��  ]rc�  (j��  ]rd�  (h	h�e]re�  (hh<e]rf�  (hhe]rg�  (j��  ]rh�  (h	h
e]ri�  (hh�e]rj�  (hhe]rk�  (j�  ]rl�  (h	h�e]rm�  (hh�eeee]rn�  (hhee]ro�  (h!]rp�  (h#h$e]rq�  (h	h�e]rr�  (hh�e]rs�  (h)heeeja�  ja�  ]rt�  (j��  ]ru�  (j��  ]rv�  (j��  ]rw�  (h	h�e]rx�  (hh<e]ry�  (hhe]rz�  (j��  ]r{�  (h	h
e]r|�  (hh�e]r}�  (hhe]r~�  (j�  ]r�  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeejt�  jt�  jt�  jt�  jt�  jt�  jt�  jt�  jt�  jt�  jt�  jt�  jt�  jt�  jt�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  ]r��  (j��  ]r��  (j��  ]r²  (j��  ]rò  (h	h�e]rĲ  (hh<e]rŲ  (hhe]rƲ  (j��  ]rǲ  (h	h
e]rȲ  (hh�e]rɲ  (hhe]rʲ  (j�  ]r˲  (h	h�e]r̲  (hh�eeee]rͲ  (hhee]rβ  (h!]rϲ  (h#h$e]rв  (h	h�e]rѲ  (hh�e]rҲ  (h)heee]rӲ  (j��  ]rԲ  (j��  ]rղ  (j��  ]rֲ  (h	h�e]rײ  (hh<e]rز  (hhe]rٲ  (j��  ]rڲ  (h	h
e]r۲  (hh�e]rܲ  (hhe]rݲ  (j�  ]r޲  (h	h�e]r߲  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejӲ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  j�  j�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r �  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r	�  (h	h�e]r
�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  ]r�  (j��  ]r �  (j��  ]r!�  (j��  ]r"�  (h	h�e]r#�  (hh<e]r$�  (hhe]r%�  (j��  ]r&�  (h	h
e]r'�  (hh�e]r(�  (hhe]r)�  (j�  ]r*�  (h	h�e]r+�  (hh�eeee]r,�  (hhee]r-�  (h!]r.�  (h#h$e]r/�  (h	h�e]r0�  (hh�e]r1�  (h)heee]r2�  (j��  ]r3�  (j��  ]r4�  (j��  ]r5�  (h	h�e]r6�  (hh<e]r7�  (hhe]r8�  (j��  ]r9�  (h	h
e]r:�  (hh�e]r;�  (hhe]r<�  (j�  ]r=�  (h	h�e]r>�  (hh�eeee]r?�  (hhee]r@�  (h!]rA�  (h#h$e]rB�  (h	h�e]rC�  (hh�e]rD�  (h)heeej2�  j2�  j2�  j2�  j2�  j2�  j2�  ]rE�  (j��  ]rF�  (j��  ]rG�  (j��  ]rH�  (h	h�e]rI�  (hh<e]rJ�  (hhe]rK�  (j��  ]rL�  (h	h
e]rM�  (hh�e]rN�  (hhe]rO�  (j�  ]rP�  (h	h�e]rQ�  (hh�eeee]rR�  (hhee]rS�  (h!]rT�  (h#h$e]rU�  (h	h�e]rV�  (hh�e]rW�  (h)heee]rX�  (j��  ]rY�  (j��  ]rZ�  (j��  ]r[�  (h	h�e]r\�  (hh<e]r]�  (hhe]r^�  (j��  ]r_�  (h	h
e]r`�  (hh<e]ra�  (hhe]rb�  (j�  ]rc�  (h	h�e]rd�  (hh�eeee]re�  (hhee]rf�  (h!]rg�  (h#h$e]rh�  (h	h�e]ri�  (hh�e]rj�  (h)heeejX�  jX�  jX�  jX�  jX�  jX�  jX�  ]rk�  (j��  ]rl�  (j��  ]rm�  (j��  ]rn�  (h	h�e]ro�  (hh<e]rp�  (hhe]rq�  (j��  ]rr�  (h	h�e]rs�  (hh<e]rt�  (hhe]ru�  (j�  ]rv�  (h	h�e]rw�  (hh�eeee]rx�  (hhee]ry�  (h!]rz�  (h#h$e]r{�  (h	h�e]r|�  (hh�e]r}�  (h)heeejk�  ]r~�  (j��  ]r�  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej~�  j~�  j~�  j~�  j~�  j~�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r³  (h	h�e]ró  (hh�eeee]rĳ  (hhee]rų  (h!]rƳ  (h#h$e]rǳ  (h	h�e]rȳ  (hh�e]rɳ  (h)heeej��  j��  j��  ]rʳ  (j��  ]r˳  (j��  ]r̳  (j��  ]rͳ  (h	h�e]rγ  (hh<e]rϳ  (hhe]rг  (j��  ]rѳ  (h	h�e]rҳ  (hh<e]rӳ  (hhe]rԳ  (j�  ]rճ  (h	h�e]rֳ  (hh�eeee]r׳  (hhee]rس  (h!]rٳ  (h#h$e]rڳ  (h	h�e]r۳  (hh�e]rܳ  (h)heeejʳ  jʳ  ]rݳ  (j��  ]r޳  (j��  ]r߳  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejݳ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r �  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r	�  (j��  ]r
�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r �  (j�  ]r!�  (h	h�e]r"�  (hh�eeee]r#�  (hhee]r$�  (h!]r%�  (h#h$e]r&�  (h	h�e]r'�  (hh�e]r(�  (h)heeej�  j�  ]r)�  (j��  ]r*�  (j��  ]r+�  (j��  ]r,�  (h	h�e]r-�  (hh<e]r.�  (hhe]r/�  (j��  ]r0�  (h	h�e]r1�  (hh<e]r2�  (hhe]r3�  (j�  ]r4�  (h	h�e]r5�  (hh�eeee]r6�  (hhee]r7�  (h!]r8�  (h#h$e]r9�  (h	h�e]r:�  (hh�e]r;�  (h)heeej)�  ]r<�  (j��  ]r=�  (j��  ]r>�  (j��  ]r?�  (h	h�e]r@�  (hh<e]rA�  (hhe]rB�  (j��  ]rC�  (h	h�e]rD�  (hh<e]rE�  (hhe]rF�  (j�  ]rG�  (h	h�e]rH�  (hh�eeee]rI�  (hhee]rJ�  (h!]rK�  (h#h$e]rL�  (h	h�e]rM�  (hh�e]rN�  (h)heee]rO�  (j��  ]rP�  (j��  ]rQ�  (j��  ]rR�  (h	h�e]rS�  (hh<e]rT�  (hhe]rU�  (j��  ]rV�  (h	h�e]rW�  (hh<e]rX�  (hhe]rY�  (j�  ]rZ�  (h	h�e]r[�  (hh�eeee]r\�  (hhee]r]�  (h!]r^�  (h#h$e]r_�  (h	h�e]r`�  (hh�e]ra�  (h)heee]rb�  (j��  ]rc�  (j��  ]rd�  (j��  ]re�  (h	h�e]rf�  (hh<e]rg�  (hhe]rh�  (j��  ]ri�  (h	h�e]rj�  (hh<e]rk�  (hhe]rl�  (j�  ]rm�  (h	h�e]rn�  (hh�eeee]ro�  (hhee]rp�  (h!]rq�  (h#h$e]rr�  (h	h�e]rs�  (hh�e]rt�  (h)heeejb�  jb�  ]ru�  (j��  ]rv�  (j��  ]rw�  (j��  ]rx�  (h	h�e]ry�  (hh<e]rz�  (hhe]r{�  (j��  ]r|�  (h	h
e]r}�  (hh<e]r~�  (hhe]r�  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeeju�  ju�  ju�  ju�  ju�  ju�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j�  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (X	   Next-Mover��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  j��  ]r´  (j��  ]rô  (j��  ]rĴ  (j��  ]rŴ  (h	h�e]rƴ  (hh<e]rǴ  (hhe]rȴ  (j��  ]rɴ  (h	h
e]rʴ  (hh<e]r˴  (hhe]r̴  (j��  ]rʹ  (h	h�e]rδ  (hh�eeee]rϴ  (hhee]rд  (h!]rѴ  (h#h$e]rҴ  (h	h�e]rӴ  (hh�e]rԴ  (h)heeej´  j´  j´  j´  j´  j´  j´  j´  j´  j´  j´  ]rմ  (j��  ]rִ  (j��  ]r״  (j��  ]rش  (h	h�e]rٴ  (hh<e]rڴ  (hhe]r۴  (j��  ]rܴ  (h	h
e]rݴ  (hh<e]r޴  (hhe]rߴ  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejմ  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h�e]r��  (hh<e]r �  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r	�  (h!]r
�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej��  j��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r �  (h)heee]r!�  (j��  ]r"�  (j��  ]r#�  (j��  ]r$�  (h	h
e]r%�  (hh<e]r&�  (hhe]r'�  (j��  ]r(�  (h	h
e]r)�  (hh<e]r*�  (hhe]r+�  (j��  ]r,�  (h	h�e]r-�  (hh�eeee]r.�  (hhee]r/�  (h!]r0�  (h#h$e]r1�  (h	h�e]r2�  (hh�e]r3�  (h)heeej!�  ]r4�  (j��  ]r5�  (j��  ]r6�  (j��  ]r7�  (h	h
e]r8�  (hh<e]r9�  (hhe]r:�  (j��  ]r;�  (h	h
e]r<�  (hh<e]r=�  (hhe]r>�  (j��  ]r?�  (h	h�e]r@�  (hh�eeee]rA�  (hhee]rB�  (h!]rC�  (h#h$e]rD�  (h	h�e]rE�  (hh�e]rF�  (h)heee]rG�  (j��  ]rH�  (j��  ]rI�  (j��  ]rJ�  (h	h
e]rK�  (hh<e]rL�  (hhe]rM�  (j��  ]rN�  (h	h
e]rO�  (hh<e]rP�  (hhe]rQ�  (j��  ]rR�  (h	h�e]rS�  (hh�eeee]rT�  (hhee]rU�  (h!]rV�  (h#h$e]rW�  (h	h�e]rX�  (hh�e]rY�  (h)heeejG�  jG�  ]rZ�  (j��  ]r[�  (j��  ]r\�  (j��  ]r]�  (h	h
e]r^�  (hh<e]r_�  (hhe]r`�  (j��  ]ra�  (h	h
e]rb�  (hh<e]rc�  (hhe]rd�  (j��  ]re�  (h	h�e]rf�  (hh�eeee]rg�  (hhee]rh�  (h!]ri�  (h#h$e]rj�  (h	h�e]rk�  (hh�e]rl�  (h)heeejZ�  jZ�  ]rm�  (j��  ]rn�  (j��  ]ro�  (j��  ]rp�  (h	h
e]rq�  (hh<e]rr�  (hhe]rs�  (j��  ]rt�  (h	h
e]ru�  (hh<e]rv�  (hhe]rw�  (j��  ]rx�  (h	h�e]ry�  (hh�eeee]rz�  (hhee]r{�  (h!]r|�  (h#h$e]r}�  (h	h�e]r~�  (hh�e]r�  (h)heeejm�  jm�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  j��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]rµ  (hhe]rõ  (j��  ]rĵ  (h	h�e]rŵ  (hh�eeee]rƵ  (hhee]rǵ  (h!]rȵ  (h#h$e]rɵ  (h	h�e]rʵ  (hh�e]r˵  (h)heeej��  j��  j��  j��  ]r̵  (j��  ]r͵  (j��  ]rε  (j��  ]rϵ  (h	h
e]rе  (hh<e]rѵ  (hhe]rҵ  (j��  ]rӵ  (h	h
e]rԵ  (hh<e]rյ  (hhe]rֵ  (j��  ]r׵  (h	h�e]rص  (hh�eeee]rٵ  (hhee]rڵ  (h!]r۵  (h#h$e]rܵ  (h	h�e]rݵ  (hh�e]r޵  (h)heeej̵  j̵  j̵  j̵  j̵  j̵  j̵  j̵  j̵  ]rߵ  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeejߵ  jߵ  jߵ  jߵ  jߵ  jߵ  jߵ  jߵ  ]r�  (j��  ]r�  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r �  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r	�  (hh�e]r
�  (hhe]r�  (j��  ]r�  (h	h
e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej�  j�  j�  j�  j�  j�  j�  j�  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h
e]r �  (hh<e]r!�  (hhe]r"�  (j��  ]r#�  (h	h�e]r$�  (hh�eeee]r%�  (hhee]r&�  (h!]r'�  (h#h$e]r(�  (h	h�e]r)�  (hh�e]r*�  (h)heeej�  j�  ]r+�  (j��  ]r,�  (j��  ]r-�  (j��  ]r.�  (h	h
e]r/�  (hh�e]r0�  (hhe]r1�  (j��  ]r2�  (h	h
e]r3�  (hh<e]r4�  (hhe]r5�  (j��  ]r6�  (h	h�e]r7�  (hh�eeee]r8�  (hhee]r9�  (h!]r:�  (h#h$e]r;�  (h	h�e]r<�  (hh�e]r=�  (h)heeej+�  j+�  j+�  j+�  j+�  j+�  ]r>�  (j��  ]r?�  (j��  ]r@�  (j��  ]rA�  (h	h
e]rB�  (hh�e]rC�  (hhe]rD�  (j��  ]rE�  (h	h
e]rF�  (hh<e]rG�  (hhe]rH�  (j��  ]rI�  (h	h�e]rJ�  (hh�eeee]rK�  (hhee]rL�  (h!]rM�  (h#h$e]rN�  (h	h�e]rO�  (hh�e]rP�  (h)heeej>�  j>�  j>�  j>�  ]rQ�  (j��  ]rR�  (j��  ]rS�  (j��  ]rT�  (h	h
e]rU�  (hh�e]rV�  (hhe]rW�  (j��  ]rX�  (h	h
e]rY�  (hh<e]rZ�  (hhe]r[�  (j��  ]r\�  (h	h�e]r]�  (hh�eeee]r^�  (hhee]r_�  (h!]r`�  (h#h$e]ra�  (h	h�e]rb�  (hh�e]rc�  (h)heeejQ�  jQ�  jQ�  jQ�  jQ�  jQ�  jQ�  jQ�  jQ�  ]rd�  (j��  ]re�  (j��  ]rf�  (j��  ]rg�  (h	h
e]rh�  (hh�e]ri�  (hhe]rj�  (j��  ]rk�  (h	h
e]rl�  (hh<e]rm�  (hhe]rn�  (j��  ]ro�  (h	h�e]rp�  (hh�eeee]rq�  (hhee]rr�  (h!]rs�  (h#h$e]rt�  (h	h�e]ru�  (hh�e]rv�  (h)heeejd�  jd�  jd�  jd�  jd�  jd�  jd�  jd�  jd�  jd�  jd�  jd�  jd�  jd�  jd�  ]rw�  (j��  ]rx�  (j��  ]ry�  (j��  ]rz�  (h	h
e]r{�  (hh�e]r|�  (hhe]r}�  (j��  ]r~�  (h	h
e]r�  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeejw�  jw�  jw�  jw�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej��  j��  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heee]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r��  (hh�e]r��  (hhe]r��  (j��  ]r��  (h	h
e]r��  (hh<e]r��  (hhe]r��  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r¶  (h)heee]rö  (j��  ]rĶ  (j��  ]rŶ  (j��  ]rƶ  (h	h
e]rǶ  (hh�e]rȶ  (hhe]rɶ  (j��  ]rʶ  (h	h
e]r˶  (hh<e]r̶  (hhe]rͶ  (j��  ]rζ  (h	h�e]r϶  (hh�eeee]rж  (hhee]rѶ  (h!]rҶ  (h#h$e]rӶ  (h	h�e]rԶ  (hh�e]rն  (h)heee]rֶ  (j��  ]r׶  (j��  ]rض  (j��  ]rٶ  (h	h
e]rڶ  (hh�e]r۶  (hhe]rܶ  (j��  ]rݶ  (h	h
e]r޶  (hh<e]r߶  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heee]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r��  (h	h�e]r��  (hh�eeee]r��  (hhee]r��  (h!]r��  (h#h$e]r��  (h	h�e]r��  (hh�e]r��  (h)heeej�  j�  j�  j�  ]r��  (j��  ]r��  (j��  ]r��  (j��  ]r��  (h	h
e]r �  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh�eeee]r	�  (hhee]r
�  (h!]r�  (h#h$e]r�  (h	h�e]r�  (hh�e]r�  (h)heeej��  ]r�  (j��  ]r�  (j��  ]r�  (j��  ]r�  (h	h
e]r�  (hh�e]r�  (hhe]r�  (j��  ]r�  (h	h�e]r�  (hh<e]r�  (hhe]r�  (X	   Next-Mover�  ]r�  (h	h�e]r�  (hh�eeee]r�  (hhee]r�  (h!]r�  (h#h$e]r �  (h	h�e]r!�  (hh�e]r"�  (h)heeej�  e(]r#�  (j��  ]r$�  (j��  ]r%�  (j��  ]r&�  (h	h
e]r'�  (hh�e]r(�  (hhe]r)�  (j��  ]r*�  (h	h�e]r+�  (hh<e]r,�  (hhe]r-�  (j�  ]r.�  (h	h�e]r/�  (hh�eeee]r0�  (hhee]r1�  (h!]r2�  (h#h$e]r3�  (h	h�e]r4�  (hh�e]r5�  (h)heeeee.