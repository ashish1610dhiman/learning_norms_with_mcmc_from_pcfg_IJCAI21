�]q (X   Normsq]q(X   Proq]q(X   Performq]q(X   ZoneqX   2qe]q	(X   Actionq
X   putdownqee]q(X   Onq]q(X   ColourqX   bqe]q(X   ShapeqX   circleqeee]q(X   Perq]q(h]q(hX   1qe]q(h
X   putdownqee]q(h]q(hX   rqe]q(hX   squareqeeee.